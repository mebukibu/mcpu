module ram (clk, load, addr, d, q);

  input clk, load;
  input [15:0] addr;
  input [7:0] d;
  output [7:0] q;
  reg [7:0] mem[0:2**16-1];

  assign q = mem[addr];

  always @(posedge clk)
    if (load)
      mem[addr] <= d;

  initial begin
    mem[16'h0000] = 8'h22; // JMP main
    mem[16'h0001] = 8'hCE;
    mem[16'h0002] = 8'h1C;
    mem[16'h0003] = 8'h00;
    mem[16'h0004] = 8'h00;
    mem[16'h0005] = 8'h00;
    mem[16'h0006] = 8'h00;
    mem[16'h0007] = 8'h00;
    mem[16'h0008] = 8'h00;
                          // pos:
    mem[16'h0009] = 8'h00;
    mem[16'h000A] = 8'h00;
    mem[16'h000B] = 8'h00;
    mem[16'h000C] = 8'h00;
    mem[16'h000D] = 8'h00;
    mem[16'h000E] = 8'h00;
    mem[16'h000F] = 8'h00;
    mem[16'h0010] = 8'h00;
    mem[16'h0011] = 8'h00;
    mem[16'h0012] = 8'h00;
    mem[16'h0013] = 8'h00;
    mem[16'h0014] = 8'h00;
    mem[16'h0015] = 8'h00;
    mem[16'h0016] = 8'h00;
    mem[16'h0017] = 8'h00;
    mem[16'h0018] = 8'h00;
    mem[16'h0019] = 8'h00;
    mem[16'h001A] = 8'h00;
    mem[16'h001B] = 8'h00;
    mem[16'h001C] = 8'h00;
    mem[16'h001D] = 8'h00;
    mem[16'h001E] = 8'h00;
    mem[16'h001F] = 8'h00;
    mem[16'h0020] = 8'h00;
    mem[16'h0021] = 8'h00;
    mem[16'h0022] = 8'h00;
    mem[16'h0023] = 8'h00;
    mem[16'h0024] = 8'h00;
    mem[16'h0025] = 8'h00;
    mem[16'h0026] = 8'h00;
    mem[16'h0027] = 8'h00;
    mem[16'h0028] = 8'h00;
    mem[16'h0029] = 8'h00;
    mem[16'h002A] = 8'h00;
    mem[16'h002B] = 8'h00;
    mem[16'h002C] = 8'h00;
    mem[16'h002D] = 8'h00;
    mem[16'h002E] = 8'h00;
    mem[16'h002F] = 8'h00;
    mem[16'h0030] = 8'h00;
    mem[16'h0031] = 8'h00;
    mem[16'h0032] = 8'h00;
    mem[16'h0033] = 8'h00;
    mem[16'h0034] = 8'h00;
    mem[16'h0035] = 8'h00;
    mem[16'h0036] = 8'h00;
    mem[16'h0037] = 8'h00;
    mem[16'h0038] = 8'h00;
    mem[16'h0039] = 8'h00;
    mem[16'h003A] = 8'h00;
    mem[16'h003B] = 8'h00;
    mem[16'h003C] = 8'h00;
    mem[16'h003D] = 8'h00;
    mem[16'h003E] = 8'h00;
    mem[16'h003F] = 8'h00;
    mem[16'h0040] = 8'h00;
    mem[16'h0041] = 8'h00;
    mem[16'h0042] = 8'h00;
    mem[16'h0043] = 8'h00;
    mem[16'h0044] = 8'h00;
    mem[16'h0045] = 8'h00;
    mem[16'h0046] = 8'h00;
    mem[16'h0047] = 8'h00;
    mem[16'h0048] = 8'h00;
                          // check:
    mem[16'h0049] = 8'h85; // SUBN RSP 8
    mem[16'h004A] = 8'h06;
    mem[16'h004B] = 8'h08;
    mem[16'h004C] = 8'h00;
    mem[16'h004D] = 8'h00;
    mem[16'h004E] = 8'h00;
    mem[16'h004F] = 8'h04; // PUSH RBP
    mem[16'h0050] = 8'h05;
    mem[16'h0051] = 8'h40; // MOV RBP RSP
    mem[16'h0052] = 8'h05;
    mem[16'h0053] = 8'h06;
    mem[16'h0054] = 8'h85; // SUBN RSP 32
    mem[16'h0055] = 8'h06;
    mem[16'h0056] = 8'h20;
    mem[16'h0057] = 8'h00;
    mem[16'h0058] = 8'h00;
    mem[16'h0059] = 8'h00;
    mem[16'h005A] = 8'h40; // MOV RBX RBP
    mem[16'h005B] = 8'h07;
    mem[16'h005C] = 8'h05;
    mem[16'h005D] = 8'h85; // SUBN RBX 32
    mem[16'h005E] = 8'h07;
    mem[16'h005F] = 8'h20;
    mem[16'h0060] = 8'h00;
    mem[16'h0061] = 8'h00;
    mem[16'h0062] = 8'h00;
    mem[16'h0063] = 8'h58; // MOVAR4 RBX RDI
    mem[16'h0064] = 8'h07;
    mem[16'h0065] = 8'h01;
    mem[16'h0066] = 8'h40; // MOV RBX RBP
    mem[16'h0067] = 8'h07;
    mem[16'h0068] = 8'h05;
    mem[16'h0069] = 8'h85; // SUBN RBX 28
    mem[16'h006A] = 8'h07;
    mem[16'h006B] = 8'h1C;
    mem[16'h006C] = 8'h00;
    mem[16'h006D] = 8'h00;
    mem[16'h006E] = 8'h00;
    mem[16'h006F] = 8'h58; // MOVAR4 RBX RSI
    mem[16'h0070] = 8'h07;
    mem[16'h0071] = 8'h02;
    mem[16'h0072] = 8'h40; // MOV RBX RBP
    mem[16'h0073] = 8'h07;
    mem[16'h0074] = 8'h05;
    mem[16'h0075] = 8'h85; // SUBN RBX 24
    mem[16'h0076] = 8'h07;
    mem[16'h0077] = 8'h18;
    mem[16'h0078] = 8'h00;
    mem[16'h0079] = 8'h00;
    mem[16'h007A] = 8'h00;
    mem[16'h007B] = 8'h58; // MOVAR4 RBX RDX
    mem[16'h007C] = 8'h07;
    mem[16'h007D] = 8'h03;
    mem[16'h007E] = 8'h40; // MOV RAX RBP
    mem[16'h007F] = 8'h00;
    mem[16'h0080] = 8'h05;
    mem[16'h0081] = 8'h85; // SUBN RAX 20
    mem[16'h0082] = 8'h00;
    mem[16'h0083] = 8'h14;
    mem[16'h0084] = 8'h00;
    mem[16'h0085] = 8'h00;
    mem[16'h0086] = 8'h00;
    mem[16'h0087] = 8'h85; // SUBN RSP 8
    mem[16'h0088] = 8'h06;
    mem[16'h0089] = 8'h08;
    mem[16'h008A] = 8'h00;
    mem[16'h008B] = 8'h00;
    mem[16'h008C] = 8'h00;
    mem[16'h008D] = 8'h04; // PUSH RAX
    mem[16'h008E] = 8'h00;
    mem[16'h008F] = 8'h85; // SUBN RSP 8
    mem[16'h0090] = 8'h06;
    mem[16'h0091] = 8'h08;
    mem[16'h0092] = 8'h00;
    mem[16'h0093] = 8'h00;
    mem[16'h0094] = 8'h00;
    mem[16'h0095] = 8'h05; // PUSHN 0
    mem[16'h0096] = 8'h00;
    mem[16'h0097] = 8'h00;
    mem[16'h0098] = 8'h00;
    mem[16'h0099] = 8'h00;
    mem[16'h009A] = 8'h00;
    mem[16'h009B] = 8'h08; // POP RDI
    mem[16'h009C] = 8'h01;
    mem[16'h009D] = 8'h81; // ADDN RSP 8
    mem[16'h009E] = 8'h06;
    mem[16'h009F] = 8'h08;
    mem[16'h00A0] = 8'h00;
    mem[16'h00A1] = 8'h00;
    mem[16'h00A2] = 8'h00;
    mem[16'h00A3] = 8'h08; // POP RAX
    mem[16'h00A4] = 8'h00;
    mem[16'h00A5] = 8'h81; // ADDN RSP 8
    mem[16'h00A6] = 8'h06;
    mem[16'h00A7] = 8'h08;
    mem[16'h00A8] = 8'h00;
    mem[16'h00A9] = 8'h00;
    mem[16'h00AA] = 8'h00;
    mem[16'h00AB] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h00AC] = 8'h00;
    mem[16'h00AD] = 8'h01;
    mem[16'h00AE] = 8'h85; // SUBN RSP 8
    mem[16'h00AF] = 8'h06;
    mem[16'h00B0] = 8'h08;
    mem[16'h00B1] = 8'h00;
    mem[16'h00B2] = 8'h00;
    mem[16'h00B3] = 8'h00;
    mem[16'h00B4] = 8'h04; // PUSH RDI
    mem[16'h00B5] = 8'h01;
    mem[16'h00B6] = 8'h81; // ADDN RSP 8
    mem[16'h00B7] = 8'h06;
    mem[16'h00B8] = 8'h08;
    mem[16'h00B9] = 8'h00;
    mem[16'h00BA] = 8'h00;
    mem[16'h00BB] = 8'h00;
                          // .Lbegin0:
    mem[16'h00BC] = 8'h40; // MOV RAX RBP
    mem[16'h00BD] = 8'h00;
    mem[16'h00BE] = 8'h05;
    mem[16'h00BF] = 8'h85; // SUBN RAX 20
    mem[16'h00C0] = 8'h00;
    mem[16'h00C1] = 8'h14;
    mem[16'h00C2] = 8'h00;
    mem[16'h00C3] = 8'h00;
    mem[16'h00C4] = 8'h00;
    mem[16'h00C5] = 8'h85; // SUBN RSP 8
    mem[16'h00C6] = 8'h06;
    mem[16'h00C7] = 8'h08;
    mem[16'h00C8] = 8'h00;
    mem[16'h00C9] = 8'h00;
    mem[16'h00CA] = 8'h00;
    mem[16'h00CB] = 8'h04; // PUSH RAX
    mem[16'h00CC] = 8'h00;
    mem[16'h00CD] = 8'h08; // POP RAX
    mem[16'h00CE] = 8'h00;
    mem[16'h00CF] = 8'h81; // ADDN RSP 8
    mem[16'h00D0] = 8'h06;
    mem[16'h00D1] = 8'h08;
    mem[16'h00D2] = 8'h00;
    mem[16'h00D3] = 8'h00;
    mem[16'h00D4] = 8'h00;
    mem[16'h00D5] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h00D6] = 8'h00;
    mem[16'h00D7] = 8'h00;
    mem[16'h00D8] = 8'h85; // SUBN RSP 8
    mem[16'h00D9] = 8'h06;
    mem[16'h00DA] = 8'h08;
    mem[16'h00DB] = 8'h00;
    mem[16'h00DC] = 8'h00;
    mem[16'h00DD] = 8'h00;
    mem[16'h00DE] = 8'h04; // PUSH RAX
    mem[16'h00DF] = 8'h00;
    mem[16'h00E0] = 8'h40; // MOV RAX RBP
    mem[16'h00E1] = 8'h00;
    mem[16'h00E2] = 8'h05;
    mem[16'h00E3] = 8'h85; // SUBN RAX 24
    mem[16'h00E4] = 8'h00;
    mem[16'h00E5] = 8'h18;
    mem[16'h00E6] = 8'h00;
    mem[16'h00E7] = 8'h00;
    mem[16'h00E8] = 8'h00;
    mem[16'h00E9] = 8'h85; // SUBN RSP 8
    mem[16'h00EA] = 8'h06;
    mem[16'h00EB] = 8'h08;
    mem[16'h00EC] = 8'h00;
    mem[16'h00ED] = 8'h00;
    mem[16'h00EE] = 8'h00;
    mem[16'h00EF] = 8'h04; // PUSH RAX
    mem[16'h00F0] = 8'h00;
    mem[16'h00F1] = 8'h08; // POP RAX
    mem[16'h00F2] = 8'h00;
    mem[16'h00F3] = 8'h81; // ADDN RSP 8
    mem[16'h00F4] = 8'h06;
    mem[16'h00F5] = 8'h08;
    mem[16'h00F6] = 8'h00;
    mem[16'h00F7] = 8'h00;
    mem[16'h00F8] = 8'h00;
    mem[16'h00F9] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h00FA] = 8'h00;
    mem[16'h00FB] = 8'h00;
    mem[16'h00FC] = 8'h85; // SUBN RSP 8
    mem[16'h00FD] = 8'h06;
    mem[16'h00FE] = 8'h08;
    mem[16'h00FF] = 8'h00;
    mem[16'h0100] = 8'h00;
    mem[16'h0101] = 8'h00;
    mem[16'h0102] = 8'h04; // PUSH RAX
    mem[16'h0103] = 8'h00;
    mem[16'h0104] = 8'h08; // POP RDI
    mem[16'h0105] = 8'h01;
    mem[16'h0106] = 8'h81; // ADDN RSP 8
    mem[16'h0107] = 8'h06;
    mem[16'h0108] = 8'h08;
    mem[16'h0109] = 8'h00;
    mem[16'h010A] = 8'h00;
    mem[16'h010B] = 8'h00;
    mem[16'h010C] = 8'h08; // POP RAX
    mem[16'h010D] = 8'h00;
    mem[16'h010E] = 8'h81; // ADDN RSP 8
    mem[16'h010F] = 8'h06;
    mem[16'h0110] = 8'h08;
    mem[16'h0111] = 8'h00;
    mem[16'h0112] = 8'h00;
    mem[16'h0113] = 8'h00;
    mem[16'h0114] = 8'h90; // CMP RAX RDI
    mem[16'h0115] = 8'h00;
    mem[16'h0116] = 8'h01;
    mem[16'h0117] = 8'h18; // SETL RAX
    mem[16'h0118] = 8'h00;
    mem[16'h0119] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h011A] = 8'h00;
    mem[16'h011B] = 8'h00;
    mem[16'h011C] = 8'h85; // SUBN RSP 8
    mem[16'h011D] = 8'h06;
    mem[16'h011E] = 8'h08;
    mem[16'h011F] = 8'h00;
    mem[16'h0120] = 8'h00;
    mem[16'h0121] = 8'h00;
    mem[16'h0122] = 8'h04; // PUSH RAX
    mem[16'h0123] = 8'h00;
    mem[16'h0124] = 8'h08; // POP RAX
    mem[16'h0125] = 8'h00;
    mem[16'h0126] = 8'h81; // ADDN RSP 8
    mem[16'h0127] = 8'h06;
    mem[16'h0128] = 8'h08;
    mem[16'h0129] = 8'h00;
    mem[16'h012A] = 8'h00;
    mem[16'h012B] = 8'h00;
    mem[16'h012C] = 8'h91; // CMPN RAX 0
    mem[16'h012D] = 8'h00;
    mem[16'h012E] = 8'h00;
    mem[16'h012F] = 8'h00;
    mem[16'h0130] = 8'h00;
    mem[16'h0131] = 8'h00;
    mem[16'h0132] = 8'h26; // JE .Lend0
    mem[16'h0133] = 8'hD9;
    mem[16'h0134] = 8'h03;
    mem[16'h0135] = 8'h00;
    mem[16'h0136] = 8'h00;
    mem[16'h0137] = 8'h00;
    mem[16'h0138] = 8'h00;
    mem[16'h0139] = 8'h00;
    mem[16'h013A] = 8'h00;
    mem[16'h013B] = 8'h85; // SUBN RSP 8
    mem[16'h013C] = 8'h06;
    mem[16'h013D] = 8'h08;
    mem[16'h013E] = 8'h00;
    mem[16'h013F] = 8'h00;
    mem[16'h0140] = 8'h00;
    mem[16'h0141] = 8'h06; // PUSHA pos
    mem[16'h0142] = 8'h09;
    mem[16'h0143] = 8'h00;
    mem[16'h0144] = 8'h00;
    mem[16'h0145] = 8'h00;
    mem[16'h0146] = 8'h00;
    mem[16'h0147] = 8'h00;
    mem[16'h0148] = 8'h00;
    mem[16'h0149] = 8'h00;
    mem[16'h014A] = 8'h40; // MOV RAX RBP
    mem[16'h014B] = 8'h00;
    mem[16'h014C] = 8'h05;
    mem[16'h014D] = 8'h85; // SUBN RAX 20
    mem[16'h014E] = 8'h00;
    mem[16'h014F] = 8'h14;
    mem[16'h0150] = 8'h00;
    mem[16'h0151] = 8'h00;
    mem[16'h0152] = 8'h00;
    mem[16'h0153] = 8'h85; // SUBN RSP 8
    mem[16'h0154] = 8'h06;
    mem[16'h0155] = 8'h08;
    mem[16'h0156] = 8'h00;
    mem[16'h0157] = 8'h00;
    mem[16'h0158] = 8'h00;
    mem[16'h0159] = 8'h04; // PUSH RAX
    mem[16'h015A] = 8'h00;
    mem[16'h015B] = 8'h08; // POP RAX
    mem[16'h015C] = 8'h00;
    mem[16'h015D] = 8'h81; // ADDN RSP 8
    mem[16'h015E] = 8'h06;
    mem[16'h015F] = 8'h08;
    mem[16'h0160] = 8'h00;
    mem[16'h0161] = 8'h00;
    mem[16'h0162] = 8'h00;
    mem[16'h0163] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0164] = 8'h00;
    mem[16'h0165] = 8'h00;
    mem[16'h0166] = 8'h85; // SUBN RSP 8
    mem[16'h0167] = 8'h06;
    mem[16'h0168] = 8'h08;
    mem[16'h0169] = 8'h00;
    mem[16'h016A] = 8'h00;
    mem[16'h016B] = 8'h00;
    mem[16'h016C] = 8'h04; // PUSH RAX
    mem[16'h016D] = 8'h00;
    mem[16'h016E] = 8'h08; // POP RDI
    mem[16'h016F] = 8'h01;
    mem[16'h0170] = 8'h81; // ADDN RSP 8
    mem[16'h0171] = 8'h06;
    mem[16'h0172] = 8'h08;
    mem[16'h0173] = 8'h00;
    mem[16'h0174] = 8'h00;
    mem[16'h0175] = 8'h00;
    mem[16'h0176] = 8'h08; // POP RAX
    mem[16'h0177] = 8'h00;
    mem[16'h0178] = 8'h81; // ADDN RSP 8
    mem[16'h0179] = 8'h06;
    mem[16'h017A] = 8'h08;
    mem[16'h017B] = 8'h00;
    mem[16'h017C] = 8'h00;
    mem[16'h017D] = 8'h00;
    mem[16'h017E] = 8'h89; // MULN RDI 8
    mem[16'h017F] = 8'h01;
    mem[16'h0180] = 8'h08;
    mem[16'h0181] = 8'h00;
    mem[16'h0182] = 8'h00;
    mem[16'h0183] = 8'h00;
    mem[16'h0184] = 8'h80; // ADD RAX RDI
    mem[16'h0185] = 8'h00;
    mem[16'h0186] = 8'h01;
    mem[16'h0187] = 8'h85; // SUBN RSP 8
    mem[16'h0188] = 8'h06;
    mem[16'h0189] = 8'h08;
    mem[16'h018A] = 8'h00;
    mem[16'h018B] = 8'h00;
    mem[16'h018C] = 8'h00;
    mem[16'h018D] = 8'h04; // PUSH RAX
    mem[16'h018E] = 8'h00;
    mem[16'h018F] = 8'h85; // SUBN RSP 8
    mem[16'h0190] = 8'h06;
    mem[16'h0191] = 8'h08;
    mem[16'h0192] = 8'h00;
    mem[16'h0193] = 8'h00;
    mem[16'h0194] = 8'h00;
    mem[16'h0195] = 8'h05; // PUSHN 0
    mem[16'h0196] = 8'h00;
    mem[16'h0197] = 8'h00;
    mem[16'h0198] = 8'h00;
    mem[16'h0199] = 8'h00;
    mem[16'h019A] = 8'h00;
    mem[16'h019B] = 8'h08; // POP RDI
    mem[16'h019C] = 8'h01;
    mem[16'h019D] = 8'h81; // ADDN RSP 8
    mem[16'h019E] = 8'h06;
    mem[16'h019F] = 8'h08;
    mem[16'h01A0] = 8'h00;
    mem[16'h01A1] = 8'h00;
    mem[16'h01A2] = 8'h00;
    mem[16'h01A3] = 8'h08; // POP RAX
    mem[16'h01A4] = 8'h00;
    mem[16'h01A5] = 8'h81; // ADDN RSP 8
    mem[16'h01A6] = 8'h06;
    mem[16'h01A7] = 8'h08;
    mem[16'h01A8] = 8'h00;
    mem[16'h01A9] = 8'h00;
    mem[16'h01AA] = 8'h00;
    mem[16'h01AB] = 8'h89; // MULN RDI 4
    mem[16'h01AC] = 8'h01;
    mem[16'h01AD] = 8'h04;
    mem[16'h01AE] = 8'h00;
    mem[16'h01AF] = 8'h00;
    mem[16'h01B0] = 8'h00;
    mem[16'h01B1] = 8'h80; // ADD RAX RDI
    mem[16'h01B2] = 8'h00;
    mem[16'h01B3] = 8'h01;
    mem[16'h01B4] = 8'h85; // SUBN RSP 8
    mem[16'h01B5] = 8'h06;
    mem[16'h01B6] = 8'h08;
    mem[16'h01B7] = 8'h00;
    mem[16'h01B8] = 8'h00;
    mem[16'h01B9] = 8'h00;
    mem[16'h01BA] = 8'h04; // PUSH RAX
    mem[16'h01BB] = 8'h00;
    mem[16'h01BC] = 8'h08; // POP RAX
    mem[16'h01BD] = 8'h00;
    mem[16'h01BE] = 8'h81; // ADDN RSP 8
    mem[16'h01BF] = 8'h06;
    mem[16'h01C0] = 8'h08;
    mem[16'h01C1] = 8'h00;
    mem[16'h01C2] = 8'h00;
    mem[16'h01C3] = 8'h00;
    mem[16'h01C4] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h01C5] = 8'h00;
    mem[16'h01C6] = 8'h00;
    mem[16'h01C7] = 8'h85; // SUBN RSP 8
    mem[16'h01C8] = 8'h06;
    mem[16'h01C9] = 8'h08;
    mem[16'h01CA] = 8'h00;
    mem[16'h01CB] = 8'h00;
    mem[16'h01CC] = 8'h00;
    mem[16'h01CD] = 8'h04; // PUSH RAX
    mem[16'h01CE] = 8'h00;
    mem[16'h01CF] = 8'h40; // MOV RAX RBP
    mem[16'h01D0] = 8'h00;
    mem[16'h01D1] = 8'h05;
    mem[16'h01D2] = 8'h85; // SUBN RAX 32
    mem[16'h01D3] = 8'h00;
    mem[16'h01D4] = 8'h20;
    mem[16'h01D5] = 8'h00;
    mem[16'h01D6] = 8'h00;
    mem[16'h01D7] = 8'h00;
    mem[16'h01D8] = 8'h85; // SUBN RSP 8
    mem[16'h01D9] = 8'h06;
    mem[16'h01DA] = 8'h08;
    mem[16'h01DB] = 8'h00;
    mem[16'h01DC] = 8'h00;
    mem[16'h01DD] = 8'h00;
    mem[16'h01DE] = 8'h04; // PUSH RAX
    mem[16'h01DF] = 8'h00;
    mem[16'h01E0] = 8'h08; // POP RAX
    mem[16'h01E1] = 8'h00;
    mem[16'h01E2] = 8'h81; // ADDN RSP 8
    mem[16'h01E3] = 8'h06;
    mem[16'h01E4] = 8'h08;
    mem[16'h01E5] = 8'h00;
    mem[16'h01E6] = 8'h00;
    mem[16'h01E7] = 8'h00;
    mem[16'h01E8] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h01E9] = 8'h00;
    mem[16'h01EA] = 8'h00;
    mem[16'h01EB] = 8'h85; // SUBN RSP 8
    mem[16'h01EC] = 8'h06;
    mem[16'h01ED] = 8'h08;
    mem[16'h01EE] = 8'h00;
    mem[16'h01EF] = 8'h00;
    mem[16'h01F0] = 8'h00;
    mem[16'h01F1] = 8'h04; // PUSH RAX
    mem[16'h01F2] = 8'h00;
    mem[16'h01F3] = 8'h08; // POP RDI
    mem[16'h01F4] = 8'h01;
    mem[16'h01F5] = 8'h81; // ADDN RSP 8
    mem[16'h01F6] = 8'h06;
    mem[16'h01F7] = 8'h08;
    mem[16'h01F8] = 8'h00;
    mem[16'h01F9] = 8'h00;
    mem[16'h01FA] = 8'h00;
    mem[16'h01FB] = 8'h08; // POP RAX
    mem[16'h01FC] = 8'h00;
    mem[16'h01FD] = 8'h81; // ADDN RSP 8
    mem[16'h01FE] = 8'h06;
    mem[16'h01FF] = 8'h08;
    mem[16'h0200] = 8'h00;
    mem[16'h0201] = 8'h00;
    mem[16'h0202] = 8'h00;
    mem[16'h0203] = 8'h90; // CMP RAX RDI
    mem[16'h0204] = 8'h00;
    mem[16'h0205] = 8'h01;
    mem[16'h0206] = 8'h10; // SETE RAX
    mem[16'h0207] = 8'h00;
    mem[16'h0208] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h0209] = 8'h00;
    mem[16'h020A] = 8'h00;
    mem[16'h020B] = 8'h85; // SUBN RSP 8
    mem[16'h020C] = 8'h06;
    mem[16'h020D] = 8'h08;
    mem[16'h020E] = 8'h00;
    mem[16'h020F] = 8'h00;
    mem[16'h0210] = 8'h00;
    mem[16'h0211] = 8'h04; // PUSH RAX
    mem[16'h0212] = 8'h00;
    mem[16'h0213] = 8'h08; // POP RAX
    mem[16'h0214] = 8'h00;
    mem[16'h0215] = 8'h81; // ADDN RSP 8
    mem[16'h0216] = 8'h06;
    mem[16'h0217] = 8'h08;
    mem[16'h0218] = 8'h00;
    mem[16'h0219] = 8'h00;
    mem[16'h021A] = 8'h00;
    mem[16'h021B] = 8'h91; // CMPN RAX 0
    mem[16'h021C] = 8'h00;
    mem[16'h021D] = 8'h00;
    mem[16'h021E] = 8'h00;
    mem[16'h021F] = 8'h00;
    mem[16'h0220] = 8'h00;
    mem[16'h0221] = 8'h26; // JE .Lend1
    mem[16'h0222] = 8'h47;
    mem[16'h0223] = 8'h02;
    mem[16'h0224] = 8'h00;
    mem[16'h0225] = 8'h00;
    mem[16'h0226] = 8'h00;
    mem[16'h0227] = 8'h00;
    mem[16'h0228] = 8'h00;
    mem[16'h0229] = 8'h00;
    mem[16'h022A] = 8'h85; // SUBN RSP 8
    mem[16'h022B] = 8'h06;
    mem[16'h022C] = 8'h08;
    mem[16'h022D] = 8'h00;
    mem[16'h022E] = 8'h00;
    mem[16'h022F] = 8'h00;
    mem[16'h0230] = 8'h05; // PUSHN 0
    mem[16'h0231] = 8'h00;
    mem[16'h0232] = 8'h00;
    mem[16'h0233] = 8'h00;
    mem[16'h0234] = 8'h00;
    mem[16'h0235] = 8'h00;
    mem[16'h0236] = 8'h08; // POP RAX
    mem[16'h0237] = 8'h00;
    mem[16'h0238] = 8'h81; // ADDN RSP 8
    mem[16'h0239] = 8'h06;
    mem[16'h023A] = 8'h08;
    mem[16'h023B] = 8'h00;
    mem[16'h023C] = 8'h00;
    mem[16'h023D] = 8'h00;
    mem[16'h023E] = 8'h22; // JMP .Lreturn.check
    mem[16'h023F] = 8'h08;
    mem[16'h0240] = 8'h16;
    mem[16'h0241] = 8'h00;
    mem[16'h0242] = 8'h00;
    mem[16'h0243] = 8'h00;
    mem[16'h0244] = 8'h00;
    mem[16'h0245] = 8'h00;
    mem[16'h0246] = 8'h00;
                          // .Lend1:
    mem[16'h0247] = 8'h85; // SUBN RSP 8
    mem[16'h0248] = 8'h06;
    mem[16'h0249] = 8'h08;
    mem[16'h024A] = 8'h00;
    mem[16'h024B] = 8'h00;
    mem[16'h024C] = 8'h00;
    mem[16'h024D] = 8'h06; // PUSHA pos
    mem[16'h024E] = 8'h09;
    mem[16'h024F] = 8'h00;
    mem[16'h0250] = 8'h00;
    mem[16'h0251] = 8'h00;
    mem[16'h0252] = 8'h00;
    mem[16'h0253] = 8'h00;
    mem[16'h0254] = 8'h00;
    mem[16'h0255] = 8'h00;
    mem[16'h0256] = 8'h40; // MOV RAX RBP
    mem[16'h0257] = 8'h00;
    mem[16'h0258] = 8'h05;
    mem[16'h0259] = 8'h85; // SUBN RAX 20
    mem[16'h025A] = 8'h00;
    mem[16'h025B] = 8'h14;
    mem[16'h025C] = 8'h00;
    mem[16'h025D] = 8'h00;
    mem[16'h025E] = 8'h00;
    mem[16'h025F] = 8'h85; // SUBN RSP 8
    mem[16'h0260] = 8'h06;
    mem[16'h0261] = 8'h08;
    mem[16'h0262] = 8'h00;
    mem[16'h0263] = 8'h00;
    mem[16'h0264] = 8'h00;
    mem[16'h0265] = 8'h04; // PUSH RAX
    mem[16'h0266] = 8'h00;
    mem[16'h0267] = 8'h08; // POP RAX
    mem[16'h0268] = 8'h00;
    mem[16'h0269] = 8'h81; // ADDN RSP 8
    mem[16'h026A] = 8'h06;
    mem[16'h026B] = 8'h08;
    mem[16'h026C] = 8'h00;
    mem[16'h026D] = 8'h00;
    mem[16'h026E] = 8'h00;
    mem[16'h026F] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0270] = 8'h00;
    mem[16'h0271] = 8'h00;
    mem[16'h0272] = 8'h85; // SUBN RSP 8
    mem[16'h0273] = 8'h06;
    mem[16'h0274] = 8'h08;
    mem[16'h0275] = 8'h00;
    mem[16'h0276] = 8'h00;
    mem[16'h0277] = 8'h00;
    mem[16'h0278] = 8'h04; // PUSH RAX
    mem[16'h0279] = 8'h00;
    mem[16'h027A] = 8'h08; // POP RDI
    mem[16'h027B] = 8'h01;
    mem[16'h027C] = 8'h81; // ADDN RSP 8
    mem[16'h027D] = 8'h06;
    mem[16'h027E] = 8'h08;
    mem[16'h027F] = 8'h00;
    mem[16'h0280] = 8'h00;
    mem[16'h0281] = 8'h00;
    mem[16'h0282] = 8'h08; // POP RAX
    mem[16'h0283] = 8'h00;
    mem[16'h0284] = 8'h81; // ADDN RSP 8
    mem[16'h0285] = 8'h06;
    mem[16'h0286] = 8'h08;
    mem[16'h0287] = 8'h00;
    mem[16'h0288] = 8'h00;
    mem[16'h0289] = 8'h00;
    mem[16'h028A] = 8'h89; // MULN RDI 8
    mem[16'h028B] = 8'h01;
    mem[16'h028C] = 8'h08;
    mem[16'h028D] = 8'h00;
    mem[16'h028E] = 8'h00;
    mem[16'h028F] = 8'h00;
    mem[16'h0290] = 8'h80; // ADD RAX RDI
    mem[16'h0291] = 8'h00;
    mem[16'h0292] = 8'h01;
    mem[16'h0293] = 8'h85; // SUBN RSP 8
    mem[16'h0294] = 8'h06;
    mem[16'h0295] = 8'h08;
    mem[16'h0296] = 8'h00;
    mem[16'h0297] = 8'h00;
    mem[16'h0298] = 8'h00;
    mem[16'h0299] = 8'h04; // PUSH RAX
    mem[16'h029A] = 8'h00;
    mem[16'h029B] = 8'h85; // SUBN RSP 8
    mem[16'h029C] = 8'h06;
    mem[16'h029D] = 8'h08;
    mem[16'h029E] = 8'h00;
    mem[16'h029F] = 8'h00;
    mem[16'h02A0] = 8'h00;
    mem[16'h02A1] = 8'h05; // PUSHN 1
    mem[16'h02A2] = 8'h00;
    mem[16'h02A3] = 8'h01;
    mem[16'h02A4] = 8'h00;
    mem[16'h02A5] = 8'h00;
    mem[16'h02A6] = 8'h00;
    mem[16'h02A7] = 8'h08; // POP RDI
    mem[16'h02A8] = 8'h01;
    mem[16'h02A9] = 8'h81; // ADDN RSP 8
    mem[16'h02AA] = 8'h06;
    mem[16'h02AB] = 8'h08;
    mem[16'h02AC] = 8'h00;
    mem[16'h02AD] = 8'h00;
    mem[16'h02AE] = 8'h00;
    mem[16'h02AF] = 8'h08; // POP RAX
    mem[16'h02B0] = 8'h00;
    mem[16'h02B1] = 8'h81; // ADDN RSP 8
    mem[16'h02B2] = 8'h06;
    mem[16'h02B3] = 8'h08;
    mem[16'h02B4] = 8'h00;
    mem[16'h02B5] = 8'h00;
    mem[16'h02B6] = 8'h00;
    mem[16'h02B7] = 8'h89; // MULN RDI 4
    mem[16'h02B8] = 8'h01;
    mem[16'h02B9] = 8'h04;
    mem[16'h02BA] = 8'h00;
    mem[16'h02BB] = 8'h00;
    mem[16'h02BC] = 8'h00;
    mem[16'h02BD] = 8'h80; // ADD RAX RDI
    mem[16'h02BE] = 8'h00;
    mem[16'h02BF] = 8'h01;
    mem[16'h02C0] = 8'h85; // SUBN RSP 8
    mem[16'h02C1] = 8'h06;
    mem[16'h02C2] = 8'h08;
    mem[16'h02C3] = 8'h00;
    mem[16'h02C4] = 8'h00;
    mem[16'h02C5] = 8'h00;
    mem[16'h02C6] = 8'h04; // PUSH RAX
    mem[16'h02C7] = 8'h00;
    mem[16'h02C8] = 8'h08; // POP RAX
    mem[16'h02C9] = 8'h00;
    mem[16'h02CA] = 8'h81; // ADDN RSP 8
    mem[16'h02CB] = 8'h06;
    mem[16'h02CC] = 8'h08;
    mem[16'h02CD] = 8'h00;
    mem[16'h02CE] = 8'h00;
    mem[16'h02CF] = 8'h00;
    mem[16'h02D0] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h02D1] = 8'h00;
    mem[16'h02D2] = 8'h00;
    mem[16'h02D3] = 8'h85; // SUBN RSP 8
    mem[16'h02D4] = 8'h06;
    mem[16'h02D5] = 8'h08;
    mem[16'h02D6] = 8'h00;
    mem[16'h02D7] = 8'h00;
    mem[16'h02D8] = 8'h00;
    mem[16'h02D9] = 8'h04; // PUSH RAX
    mem[16'h02DA] = 8'h00;
    mem[16'h02DB] = 8'h40; // MOV RAX RBP
    mem[16'h02DC] = 8'h00;
    mem[16'h02DD] = 8'h05;
    mem[16'h02DE] = 8'h85; // SUBN RAX 28
    mem[16'h02DF] = 8'h00;
    mem[16'h02E0] = 8'h1C;
    mem[16'h02E1] = 8'h00;
    mem[16'h02E2] = 8'h00;
    mem[16'h02E3] = 8'h00;
    mem[16'h02E4] = 8'h85; // SUBN RSP 8
    mem[16'h02E5] = 8'h06;
    mem[16'h02E6] = 8'h08;
    mem[16'h02E7] = 8'h00;
    mem[16'h02E8] = 8'h00;
    mem[16'h02E9] = 8'h00;
    mem[16'h02EA] = 8'h04; // PUSH RAX
    mem[16'h02EB] = 8'h00;
    mem[16'h02EC] = 8'h08; // POP RAX
    mem[16'h02ED] = 8'h00;
    mem[16'h02EE] = 8'h81; // ADDN RSP 8
    mem[16'h02EF] = 8'h06;
    mem[16'h02F0] = 8'h08;
    mem[16'h02F1] = 8'h00;
    mem[16'h02F2] = 8'h00;
    mem[16'h02F3] = 8'h00;
    mem[16'h02F4] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h02F5] = 8'h00;
    mem[16'h02F6] = 8'h00;
    mem[16'h02F7] = 8'h85; // SUBN RSP 8
    mem[16'h02F8] = 8'h06;
    mem[16'h02F9] = 8'h08;
    mem[16'h02FA] = 8'h00;
    mem[16'h02FB] = 8'h00;
    mem[16'h02FC] = 8'h00;
    mem[16'h02FD] = 8'h04; // PUSH RAX
    mem[16'h02FE] = 8'h00;
    mem[16'h02FF] = 8'h08; // POP RDI
    mem[16'h0300] = 8'h01;
    mem[16'h0301] = 8'h81; // ADDN RSP 8
    mem[16'h0302] = 8'h06;
    mem[16'h0303] = 8'h08;
    mem[16'h0304] = 8'h00;
    mem[16'h0305] = 8'h00;
    mem[16'h0306] = 8'h00;
    mem[16'h0307] = 8'h08; // POP RAX
    mem[16'h0308] = 8'h00;
    mem[16'h0309] = 8'h81; // ADDN RSP 8
    mem[16'h030A] = 8'h06;
    mem[16'h030B] = 8'h08;
    mem[16'h030C] = 8'h00;
    mem[16'h030D] = 8'h00;
    mem[16'h030E] = 8'h00;
    mem[16'h030F] = 8'h90; // CMP RAX RDI
    mem[16'h0310] = 8'h00;
    mem[16'h0311] = 8'h01;
    mem[16'h0312] = 8'h10; // SETE RAX
    mem[16'h0313] = 8'h00;
    mem[16'h0314] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h0315] = 8'h00;
    mem[16'h0316] = 8'h00;
    mem[16'h0317] = 8'h85; // SUBN RSP 8
    mem[16'h0318] = 8'h06;
    mem[16'h0319] = 8'h08;
    mem[16'h031A] = 8'h00;
    mem[16'h031B] = 8'h00;
    mem[16'h031C] = 8'h00;
    mem[16'h031D] = 8'h04; // PUSH RAX
    mem[16'h031E] = 8'h00;
    mem[16'h031F] = 8'h08; // POP RAX
    mem[16'h0320] = 8'h00;
    mem[16'h0321] = 8'h81; // ADDN RSP 8
    mem[16'h0322] = 8'h06;
    mem[16'h0323] = 8'h08;
    mem[16'h0324] = 8'h00;
    mem[16'h0325] = 8'h00;
    mem[16'h0326] = 8'h00;
    mem[16'h0327] = 8'h91; // CMPN RAX 0
    mem[16'h0328] = 8'h00;
    mem[16'h0329] = 8'h00;
    mem[16'h032A] = 8'h00;
    mem[16'h032B] = 8'h00;
    mem[16'h032C] = 8'h00;
    mem[16'h032D] = 8'h26; // JE .Lend2
    mem[16'h032E] = 8'h53;
    mem[16'h032F] = 8'h03;
    mem[16'h0330] = 8'h00;
    mem[16'h0331] = 8'h00;
    mem[16'h0332] = 8'h00;
    mem[16'h0333] = 8'h00;
    mem[16'h0334] = 8'h00;
    mem[16'h0335] = 8'h00;
    mem[16'h0336] = 8'h85; // SUBN RSP 8
    mem[16'h0337] = 8'h06;
    mem[16'h0338] = 8'h08;
    mem[16'h0339] = 8'h00;
    mem[16'h033A] = 8'h00;
    mem[16'h033B] = 8'h00;
    mem[16'h033C] = 8'h05; // PUSHN 0
    mem[16'h033D] = 8'h00;
    mem[16'h033E] = 8'h00;
    mem[16'h033F] = 8'h00;
    mem[16'h0340] = 8'h00;
    mem[16'h0341] = 8'h00;
    mem[16'h0342] = 8'h08; // POP RAX
    mem[16'h0343] = 8'h00;
    mem[16'h0344] = 8'h81; // ADDN RSP 8
    mem[16'h0345] = 8'h06;
    mem[16'h0346] = 8'h08;
    mem[16'h0347] = 8'h00;
    mem[16'h0348] = 8'h00;
    mem[16'h0349] = 8'h00;
    mem[16'h034A] = 8'h22; // JMP .Lreturn.check
    mem[16'h034B] = 8'h08;
    mem[16'h034C] = 8'h16;
    mem[16'h034D] = 8'h00;
    mem[16'h034E] = 8'h00;
    mem[16'h034F] = 8'h00;
    mem[16'h0350] = 8'h00;
    mem[16'h0351] = 8'h00;
    mem[16'h0352] = 8'h00;
                          // .Lend2:
    mem[16'h0353] = 8'h40; // MOV RAX RBP
    mem[16'h0354] = 8'h00;
    mem[16'h0355] = 8'h05;
    mem[16'h0356] = 8'h85; // SUBN RAX 20
    mem[16'h0357] = 8'h00;
    mem[16'h0358] = 8'h14;
    mem[16'h0359] = 8'h00;
    mem[16'h035A] = 8'h00;
    mem[16'h035B] = 8'h00;
    mem[16'h035C] = 8'h85; // SUBN RSP 8
    mem[16'h035D] = 8'h06;
    mem[16'h035E] = 8'h08;
    mem[16'h035F] = 8'h00;
    mem[16'h0360] = 8'h00;
    mem[16'h0361] = 8'h00;
    mem[16'h0362] = 8'h04; // PUSH RAX
    mem[16'h0363] = 8'h00;
    mem[16'h0364] = 8'h40; // MOV RAX RBP
    mem[16'h0365] = 8'h00;
    mem[16'h0366] = 8'h05;
    mem[16'h0367] = 8'h85; // SUBN RAX 20
    mem[16'h0368] = 8'h00;
    mem[16'h0369] = 8'h14;
    mem[16'h036A] = 8'h00;
    mem[16'h036B] = 8'h00;
    mem[16'h036C] = 8'h00;
    mem[16'h036D] = 8'h85; // SUBN RSP 8
    mem[16'h036E] = 8'h06;
    mem[16'h036F] = 8'h08;
    mem[16'h0370] = 8'h00;
    mem[16'h0371] = 8'h00;
    mem[16'h0372] = 8'h00;
    mem[16'h0373] = 8'h04; // PUSH RAX
    mem[16'h0374] = 8'h00;
    mem[16'h0375] = 8'h08; // POP RAX
    mem[16'h0376] = 8'h00;
    mem[16'h0377] = 8'h81; // ADDN RSP 8
    mem[16'h0378] = 8'h06;
    mem[16'h0379] = 8'h08;
    mem[16'h037A] = 8'h00;
    mem[16'h037B] = 8'h00;
    mem[16'h037C] = 8'h00;
    mem[16'h037D] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h037E] = 8'h00;
    mem[16'h037F] = 8'h00;
    mem[16'h0380] = 8'h85; // SUBN RSP 8
    mem[16'h0381] = 8'h06;
    mem[16'h0382] = 8'h08;
    mem[16'h0383] = 8'h00;
    mem[16'h0384] = 8'h00;
    mem[16'h0385] = 8'h00;
    mem[16'h0386] = 8'h04; // PUSH RAX
    mem[16'h0387] = 8'h00;
    mem[16'h0388] = 8'h85; // SUBN RSP 8
    mem[16'h0389] = 8'h06;
    mem[16'h038A] = 8'h08;
    mem[16'h038B] = 8'h00;
    mem[16'h038C] = 8'h00;
    mem[16'h038D] = 8'h00;
    mem[16'h038E] = 8'h05; // PUSHN 1
    mem[16'h038F] = 8'h00;
    mem[16'h0390] = 8'h01;
    mem[16'h0391] = 8'h00;
    mem[16'h0392] = 8'h00;
    mem[16'h0393] = 8'h00;
    mem[16'h0394] = 8'h08; // POP RDI
    mem[16'h0395] = 8'h01;
    mem[16'h0396] = 8'h81; // ADDN RSP 8
    mem[16'h0397] = 8'h06;
    mem[16'h0398] = 8'h08;
    mem[16'h0399] = 8'h00;
    mem[16'h039A] = 8'h00;
    mem[16'h039B] = 8'h00;
    mem[16'h039C] = 8'h08; // POP RAX
    mem[16'h039D] = 8'h00;
    mem[16'h039E] = 8'h81; // ADDN RSP 8
    mem[16'h039F] = 8'h06;
    mem[16'h03A0] = 8'h08;
    mem[16'h03A1] = 8'h00;
    mem[16'h03A2] = 8'h00;
    mem[16'h03A3] = 8'h00;
    mem[16'h03A4] = 8'h80; // ADD RAX RDI
    mem[16'h03A5] = 8'h00;
    mem[16'h03A6] = 8'h01;
    mem[16'h03A7] = 8'h85; // SUBN RSP 8
    mem[16'h03A8] = 8'h06;
    mem[16'h03A9] = 8'h08;
    mem[16'h03AA] = 8'h00;
    mem[16'h03AB] = 8'h00;
    mem[16'h03AC] = 8'h00;
    mem[16'h03AD] = 8'h04; // PUSH RAX
    mem[16'h03AE] = 8'h00;
    mem[16'h03AF] = 8'h08; // POP RDI
    mem[16'h03B0] = 8'h01;
    mem[16'h03B1] = 8'h81; // ADDN RSP 8
    mem[16'h03B2] = 8'h06;
    mem[16'h03B3] = 8'h08;
    mem[16'h03B4] = 8'h00;
    mem[16'h03B5] = 8'h00;
    mem[16'h03B6] = 8'h00;
    mem[16'h03B7] = 8'h08; // POP RAX
    mem[16'h03B8] = 8'h00;
    mem[16'h03B9] = 8'h81; // ADDN RSP 8
    mem[16'h03BA] = 8'h06;
    mem[16'h03BB] = 8'h08;
    mem[16'h03BC] = 8'h00;
    mem[16'h03BD] = 8'h00;
    mem[16'h03BE] = 8'h00;
    mem[16'h03BF] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h03C0] = 8'h00;
    mem[16'h03C1] = 8'h01;
    mem[16'h03C2] = 8'h85; // SUBN RSP 8
    mem[16'h03C3] = 8'h06;
    mem[16'h03C4] = 8'h08;
    mem[16'h03C5] = 8'h00;
    mem[16'h03C6] = 8'h00;
    mem[16'h03C7] = 8'h00;
    mem[16'h03C8] = 8'h04; // PUSH RDI
    mem[16'h03C9] = 8'h01;
    mem[16'h03CA] = 8'h81; // ADDN RSP 8
    mem[16'h03CB] = 8'h06;
    mem[16'h03CC] = 8'h08;
    mem[16'h03CD] = 8'h00;
    mem[16'h03CE] = 8'h00;
    mem[16'h03CF] = 8'h00;
    mem[16'h03D0] = 8'h22; // JMP .Lbegin0
    mem[16'h03D1] = 8'hBC;
    mem[16'h03D2] = 8'h00;
    mem[16'h03D3] = 8'h00;
    mem[16'h03D4] = 8'h00;
    mem[16'h03D5] = 8'h00;
    mem[16'h03D6] = 8'h00;
    mem[16'h03D7] = 8'h00;
    mem[16'h03D8] = 8'h00;
                          // .Lend0:
    mem[16'h03D9] = 8'h40; // MOV RAX RBP
    mem[16'h03DA] = 8'h00;
    mem[16'h03DB] = 8'h05;
    mem[16'h03DC] = 8'h85; // SUBN RAX 28
    mem[16'h03DD] = 8'h00;
    mem[16'h03DE] = 8'h1C;
    mem[16'h03DF] = 8'h00;
    mem[16'h03E0] = 8'h00;
    mem[16'h03E1] = 8'h00;
    mem[16'h03E2] = 8'h85; // SUBN RSP 8
    mem[16'h03E3] = 8'h06;
    mem[16'h03E4] = 8'h08;
    mem[16'h03E5] = 8'h00;
    mem[16'h03E6] = 8'h00;
    mem[16'h03E7] = 8'h00;
    mem[16'h03E8] = 8'h04; // PUSH RAX
    mem[16'h03E9] = 8'h00;
    mem[16'h03EA] = 8'h08; // POP RAX
    mem[16'h03EB] = 8'h00;
    mem[16'h03EC] = 8'h81; // ADDN RSP 8
    mem[16'h03ED] = 8'h06;
    mem[16'h03EE] = 8'h08;
    mem[16'h03EF] = 8'h00;
    mem[16'h03F0] = 8'h00;
    mem[16'h03F1] = 8'h00;
    mem[16'h03F2] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h03F3] = 8'h00;
    mem[16'h03F4] = 8'h00;
    mem[16'h03F5] = 8'h85; // SUBN RSP 8
    mem[16'h03F6] = 8'h06;
    mem[16'h03F7] = 8'h08;
    mem[16'h03F8] = 8'h00;
    mem[16'h03F9] = 8'h00;
    mem[16'h03FA] = 8'h00;
    mem[16'h03FB] = 8'h04; // PUSH RAX
    mem[16'h03FC] = 8'h00;
    mem[16'h03FD] = 8'h40; // MOV RAX RBP
    mem[16'h03FE] = 8'h00;
    mem[16'h03FF] = 8'h05;
    mem[16'h0400] = 8'h85; // SUBN RAX 32
    mem[16'h0401] = 8'h00;
    mem[16'h0402] = 8'h20;
    mem[16'h0403] = 8'h00;
    mem[16'h0404] = 8'h00;
    mem[16'h0405] = 8'h00;
    mem[16'h0406] = 8'h85; // SUBN RSP 8
    mem[16'h0407] = 8'h06;
    mem[16'h0408] = 8'h08;
    mem[16'h0409] = 8'h00;
    mem[16'h040A] = 8'h00;
    mem[16'h040B] = 8'h00;
    mem[16'h040C] = 8'h04; // PUSH RAX
    mem[16'h040D] = 8'h00;
    mem[16'h040E] = 8'h08; // POP RAX
    mem[16'h040F] = 8'h00;
    mem[16'h0410] = 8'h81; // ADDN RSP 8
    mem[16'h0411] = 8'h06;
    mem[16'h0412] = 8'h08;
    mem[16'h0413] = 8'h00;
    mem[16'h0414] = 8'h00;
    mem[16'h0415] = 8'h00;
    mem[16'h0416] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0417] = 8'h00;
    mem[16'h0418] = 8'h00;
    mem[16'h0419] = 8'h85; // SUBN RSP 8
    mem[16'h041A] = 8'h06;
    mem[16'h041B] = 8'h08;
    mem[16'h041C] = 8'h00;
    mem[16'h041D] = 8'h00;
    mem[16'h041E] = 8'h00;
    mem[16'h041F] = 8'h04; // PUSH RAX
    mem[16'h0420] = 8'h00;
    mem[16'h0421] = 8'h08; // POP RDI
    mem[16'h0422] = 8'h01;
    mem[16'h0423] = 8'h81; // ADDN RSP 8
    mem[16'h0424] = 8'h06;
    mem[16'h0425] = 8'h08;
    mem[16'h0426] = 8'h00;
    mem[16'h0427] = 8'h00;
    mem[16'h0428] = 8'h00;
    mem[16'h0429] = 8'h08; // POP RAX
    mem[16'h042A] = 8'h00;
    mem[16'h042B] = 8'h81; // ADDN RSP 8
    mem[16'h042C] = 8'h06;
    mem[16'h042D] = 8'h08;
    mem[16'h042E] = 8'h00;
    mem[16'h042F] = 8'h00;
    mem[16'h0430] = 8'h00;
    mem[16'h0431] = 8'h90; // CMP RAX RDI
    mem[16'h0432] = 8'h00;
    mem[16'h0433] = 8'h01;
    mem[16'h0434] = 8'h18; // SETL RAX
    mem[16'h0435] = 8'h00;
    mem[16'h0436] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h0437] = 8'h00;
    mem[16'h0438] = 8'h00;
    mem[16'h0439] = 8'h85; // SUBN RSP 8
    mem[16'h043A] = 8'h06;
    mem[16'h043B] = 8'h08;
    mem[16'h043C] = 8'h00;
    mem[16'h043D] = 8'h00;
    mem[16'h043E] = 8'h00;
    mem[16'h043F] = 8'h04; // PUSH RAX
    mem[16'h0440] = 8'h00;
    mem[16'h0441] = 8'h08; // POP RAX
    mem[16'h0442] = 8'h00;
    mem[16'h0443] = 8'h81; // ADDN RSP 8
    mem[16'h0444] = 8'h06;
    mem[16'h0445] = 8'h08;
    mem[16'h0446] = 8'h00;
    mem[16'h0447] = 8'h00;
    mem[16'h0448] = 8'h00;
    mem[16'h0449] = 8'h91; // CMPN RAX 0
    mem[16'h044A] = 8'h00;
    mem[16'h044B] = 8'h00;
    mem[16'h044C] = 8'h00;
    mem[16'h044D] = 8'h00;
    mem[16'h044E] = 8'h00;
    mem[16'h044F] = 8'h26; // JE .Lelse3
    mem[16'h0450] = 8'hB1;
    mem[16'h0451] = 8'h05;
    mem[16'h0452] = 8'h00;
    mem[16'h0453] = 8'h00;
    mem[16'h0454] = 8'h00;
    mem[16'h0455] = 8'h00;
    mem[16'h0456] = 8'h00;
    mem[16'h0457] = 8'h00;
    mem[16'h0458] = 8'h40; // MOV RAX RBP
    mem[16'h0459] = 8'h00;
    mem[16'h045A] = 8'h05;
    mem[16'h045B] = 8'h85; // SUBN RAX 16
    mem[16'h045C] = 8'h00;
    mem[16'h045D] = 8'h10;
    mem[16'h045E] = 8'h00;
    mem[16'h045F] = 8'h00;
    mem[16'h0460] = 8'h00;
    mem[16'h0461] = 8'h85; // SUBN RSP 8
    mem[16'h0462] = 8'h06;
    mem[16'h0463] = 8'h08;
    mem[16'h0464] = 8'h00;
    mem[16'h0465] = 8'h00;
    mem[16'h0466] = 8'h00;
    mem[16'h0467] = 8'h04; // PUSH RAX
    mem[16'h0468] = 8'h00;
    mem[16'h0469] = 8'h40; // MOV RAX RBP
    mem[16'h046A] = 8'h00;
    mem[16'h046B] = 8'h05;
    mem[16'h046C] = 8'h85; // SUBN RAX 32
    mem[16'h046D] = 8'h00;
    mem[16'h046E] = 8'h20;
    mem[16'h046F] = 8'h00;
    mem[16'h0470] = 8'h00;
    mem[16'h0471] = 8'h00;
    mem[16'h0472] = 8'h85; // SUBN RSP 8
    mem[16'h0473] = 8'h06;
    mem[16'h0474] = 8'h08;
    mem[16'h0475] = 8'h00;
    mem[16'h0476] = 8'h00;
    mem[16'h0477] = 8'h00;
    mem[16'h0478] = 8'h04; // PUSH RAX
    mem[16'h0479] = 8'h00;
    mem[16'h047A] = 8'h08; // POP RAX
    mem[16'h047B] = 8'h00;
    mem[16'h047C] = 8'h81; // ADDN RSP 8
    mem[16'h047D] = 8'h06;
    mem[16'h047E] = 8'h08;
    mem[16'h047F] = 8'h00;
    mem[16'h0480] = 8'h00;
    mem[16'h0481] = 8'h00;
    mem[16'h0482] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0483] = 8'h00;
    mem[16'h0484] = 8'h00;
    mem[16'h0485] = 8'h85; // SUBN RSP 8
    mem[16'h0486] = 8'h06;
    mem[16'h0487] = 8'h08;
    mem[16'h0488] = 8'h00;
    mem[16'h0489] = 8'h00;
    mem[16'h048A] = 8'h00;
    mem[16'h048B] = 8'h04; // PUSH RAX
    mem[16'h048C] = 8'h00;
    mem[16'h048D] = 8'h40; // MOV RAX RBP
    mem[16'h048E] = 8'h00;
    mem[16'h048F] = 8'h05;
    mem[16'h0490] = 8'h85; // SUBN RAX 28
    mem[16'h0491] = 8'h00;
    mem[16'h0492] = 8'h1C;
    mem[16'h0493] = 8'h00;
    mem[16'h0494] = 8'h00;
    mem[16'h0495] = 8'h00;
    mem[16'h0496] = 8'h85; // SUBN RSP 8
    mem[16'h0497] = 8'h06;
    mem[16'h0498] = 8'h08;
    mem[16'h0499] = 8'h00;
    mem[16'h049A] = 8'h00;
    mem[16'h049B] = 8'h00;
    mem[16'h049C] = 8'h04; // PUSH RAX
    mem[16'h049D] = 8'h00;
    mem[16'h049E] = 8'h08; // POP RAX
    mem[16'h049F] = 8'h00;
    mem[16'h04A0] = 8'h81; // ADDN RSP 8
    mem[16'h04A1] = 8'h06;
    mem[16'h04A2] = 8'h08;
    mem[16'h04A3] = 8'h00;
    mem[16'h04A4] = 8'h00;
    mem[16'h04A5] = 8'h00;
    mem[16'h04A6] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h04A7] = 8'h00;
    mem[16'h04A8] = 8'h00;
    mem[16'h04A9] = 8'h85; // SUBN RSP 8
    mem[16'h04AA] = 8'h06;
    mem[16'h04AB] = 8'h08;
    mem[16'h04AC] = 8'h00;
    mem[16'h04AD] = 8'h00;
    mem[16'h04AE] = 8'h00;
    mem[16'h04AF] = 8'h04; // PUSH RAX
    mem[16'h04B0] = 8'h00;
    mem[16'h04B1] = 8'h08; // POP RDI
    mem[16'h04B2] = 8'h01;
    mem[16'h04B3] = 8'h81; // ADDN RSP 8
    mem[16'h04B4] = 8'h06;
    mem[16'h04B5] = 8'h08;
    mem[16'h04B6] = 8'h00;
    mem[16'h04B7] = 8'h00;
    mem[16'h04B8] = 8'h00;
    mem[16'h04B9] = 8'h08; // POP RAX
    mem[16'h04BA] = 8'h00;
    mem[16'h04BB] = 8'h81; // ADDN RSP 8
    mem[16'h04BC] = 8'h06;
    mem[16'h04BD] = 8'h08;
    mem[16'h04BE] = 8'h00;
    mem[16'h04BF] = 8'h00;
    mem[16'h04C0] = 8'h00;
    mem[16'h04C1] = 8'h84; // SUB RAX RDI
    mem[16'h04C2] = 8'h00;
    mem[16'h04C3] = 8'h01;
    mem[16'h04C4] = 8'h85; // SUBN RSP 8
    mem[16'h04C5] = 8'h06;
    mem[16'h04C6] = 8'h08;
    mem[16'h04C7] = 8'h00;
    mem[16'h04C8] = 8'h00;
    mem[16'h04C9] = 8'h00;
    mem[16'h04CA] = 8'h04; // PUSH RAX
    mem[16'h04CB] = 8'h00;
    mem[16'h04CC] = 8'h08; // POP RDI
    mem[16'h04CD] = 8'h01;
    mem[16'h04CE] = 8'h81; // ADDN RSP 8
    mem[16'h04CF] = 8'h06;
    mem[16'h04D0] = 8'h08;
    mem[16'h04D1] = 8'h00;
    mem[16'h04D2] = 8'h00;
    mem[16'h04D3] = 8'h00;
    mem[16'h04D4] = 8'h08; // POP RAX
    mem[16'h04D5] = 8'h00;
    mem[16'h04D6] = 8'h81; // ADDN RSP 8
    mem[16'h04D7] = 8'h06;
    mem[16'h04D8] = 8'h08;
    mem[16'h04D9] = 8'h00;
    mem[16'h04DA] = 8'h00;
    mem[16'h04DB] = 8'h00;
    mem[16'h04DC] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h04DD] = 8'h00;
    mem[16'h04DE] = 8'h01;
    mem[16'h04DF] = 8'h85; // SUBN RSP 8
    mem[16'h04E0] = 8'h06;
    mem[16'h04E1] = 8'h08;
    mem[16'h04E2] = 8'h00;
    mem[16'h04E3] = 8'h00;
    mem[16'h04E4] = 8'h00;
    mem[16'h04E5] = 8'h04; // PUSH RDI
    mem[16'h04E6] = 8'h01;
    mem[16'h04E7] = 8'h81; // ADDN RSP 8
    mem[16'h04E8] = 8'h06;
    mem[16'h04E9] = 8'h08;
    mem[16'h04EA] = 8'h00;
    mem[16'h04EB] = 8'h00;
    mem[16'h04EC] = 8'h00;
    mem[16'h04ED] = 8'h40; // MOV RAX RBP
    mem[16'h04EE] = 8'h00;
    mem[16'h04EF] = 8'h05;
    mem[16'h04F0] = 8'h85; // SUBN RAX 12
    mem[16'h04F1] = 8'h00;
    mem[16'h04F2] = 8'h0C;
    mem[16'h04F3] = 8'h00;
    mem[16'h04F4] = 8'h00;
    mem[16'h04F5] = 8'h00;
    mem[16'h04F6] = 8'h85; // SUBN RSP 8
    mem[16'h04F7] = 8'h06;
    mem[16'h04F8] = 8'h08;
    mem[16'h04F9] = 8'h00;
    mem[16'h04FA] = 8'h00;
    mem[16'h04FB] = 8'h00;
    mem[16'h04FC] = 8'h04; // PUSH RAX
    mem[16'h04FD] = 8'h00;
    mem[16'h04FE] = 8'h85; // SUBN RSP 8
    mem[16'h04FF] = 8'h06;
    mem[16'h0500] = 8'h08;
    mem[16'h0501] = 8'h00;
    mem[16'h0502] = 8'h00;
    mem[16'h0503] = 8'h00;
    mem[16'h0504] = 8'h05; // PUSHN 0
    mem[16'h0505] = 8'h00;
    mem[16'h0506] = 8'h00;
    mem[16'h0507] = 8'h00;
    mem[16'h0508] = 8'h00;
    mem[16'h0509] = 8'h00;
    mem[16'h050A] = 8'h08; // POP RDI
    mem[16'h050B] = 8'h01;
    mem[16'h050C] = 8'h81; // ADDN RSP 8
    mem[16'h050D] = 8'h06;
    mem[16'h050E] = 8'h08;
    mem[16'h050F] = 8'h00;
    mem[16'h0510] = 8'h00;
    mem[16'h0511] = 8'h00;
    mem[16'h0512] = 8'h08; // POP RAX
    mem[16'h0513] = 8'h00;
    mem[16'h0514] = 8'h81; // ADDN RSP 8
    mem[16'h0515] = 8'h06;
    mem[16'h0516] = 8'h08;
    mem[16'h0517] = 8'h00;
    mem[16'h0518] = 8'h00;
    mem[16'h0519] = 8'h00;
    mem[16'h051A] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h051B] = 8'h00;
    mem[16'h051C] = 8'h01;
    mem[16'h051D] = 8'h85; // SUBN RSP 8
    mem[16'h051E] = 8'h06;
    mem[16'h051F] = 8'h08;
    mem[16'h0520] = 8'h00;
    mem[16'h0521] = 8'h00;
    mem[16'h0522] = 8'h00;
    mem[16'h0523] = 8'h04; // PUSH RDI
    mem[16'h0524] = 8'h01;
    mem[16'h0525] = 8'h81; // ADDN RSP 8
    mem[16'h0526] = 8'h06;
    mem[16'h0527] = 8'h08;
    mem[16'h0528] = 8'h00;
    mem[16'h0529] = 8'h00;
    mem[16'h052A] = 8'h00;
    mem[16'h052B] = 8'h40; // MOV RAX RBP
    mem[16'h052C] = 8'h00;
    mem[16'h052D] = 8'h05;
    mem[16'h052E] = 8'h85; // SUBN RAX 8
    mem[16'h052F] = 8'h00;
    mem[16'h0530] = 8'h08;
    mem[16'h0531] = 8'h00;
    mem[16'h0532] = 8'h00;
    mem[16'h0533] = 8'h00;
    mem[16'h0534] = 8'h85; // SUBN RSP 8
    mem[16'h0535] = 8'h06;
    mem[16'h0536] = 8'h08;
    mem[16'h0537] = 8'h00;
    mem[16'h0538] = 8'h00;
    mem[16'h0539] = 8'h00;
    mem[16'h053A] = 8'h04; // PUSH RAX
    mem[16'h053B] = 8'h00;
    mem[16'h053C] = 8'h85; // SUBN RSP 8
    mem[16'h053D] = 8'h06;
    mem[16'h053E] = 8'h08;
    mem[16'h053F] = 8'h00;
    mem[16'h0540] = 8'h00;
    mem[16'h0541] = 8'h00;
    mem[16'h0542] = 8'h05; // PUSHN 8
    mem[16'h0543] = 8'h00;
    mem[16'h0544] = 8'h08;
    mem[16'h0545] = 8'h00;
    mem[16'h0546] = 8'h00;
    mem[16'h0547] = 8'h00;
    mem[16'h0548] = 8'h40; // MOV RAX RBP
    mem[16'h0549] = 8'h00;
    mem[16'h054A] = 8'h05;
    mem[16'h054B] = 8'h85; // SUBN RAX 16
    mem[16'h054C] = 8'h00;
    mem[16'h054D] = 8'h10;
    mem[16'h054E] = 8'h00;
    mem[16'h054F] = 8'h00;
    mem[16'h0550] = 8'h00;
    mem[16'h0551] = 8'h85; // SUBN RSP 8
    mem[16'h0552] = 8'h06;
    mem[16'h0553] = 8'h08;
    mem[16'h0554] = 8'h00;
    mem[16'h0555] = 8'h00;
    mem[16'h0556] = 8'h00;
    mem[16'h0557] = 8'h04; // PUSH RAX
    mem[16'h0558] = 8'h00;
    mem[16'h0559] = 8'h08; // POP RAX
    mem[16'h055A] = 8'h00;
    mem[16'h055B] = 8'h81; // ADDN RSP 8
    mem[16'h055C] = 8'h06;
    mem[16'h055D] = 8'h08;
    mem[16'h055E] = 8'h00;
    mem[16'h055F] = 8'h00;
    mem[16'h0560] = 8'h00;
    mem[16'h0561] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0562] = 8'h00;
    mem[16'h0563] = 8'h00;
    mem[16'h0564] = 8'h85; // SUBN RSP 8
    mem[16'h0565] = 8'h06;
    mem[16'h0566] = 8'h08;
    mem[16'h0567] = 8'h00;
    mem[16'h0568] = 8'h00;
    mem[16'h0569] = 8'h00;
    mem[16'h056A] = 8'h04; // PUSH RAX
    mem[16'h056B] = 8'h00;
    mem[16'h056C] = 8'h08; // POP RDI
    mem[16'h056D] = 8'h01;
    mem[16'h056E] = 8'h81; // ADDN RSP 8
    mem[16'h056F] = 8'h06;
    mem[16'h0570] = 8'h08;
    mem[16'h0571] = 8'h00;
    mem[16'h0572] = 8'h00;
    mem[16'h0573] = 8'h00;
    mem[16'h0574] = 8'h08; // POP RAX
    mem[16'h0575] = 8'h00;
    mem[16'h0576] = 8'h81; // ADDN RSP 8
    mem[16'h0577] = 8'h06;
    mem[16'h0578] = 8'h08;
    mem[16'h0579] = 8'h00;
    mem[16'h057A] = 8'h00;
    mem[16'h057B] = 8'h00;
    mem[16'h057C] = 8'h84; // SUB RAX RDI
    mem[16'h057D] = 8'h00;
    mem[16'h057E] = 8'h01;
    mem[16'h057F] = 8'h85; // SUBN RSP 8
    mem[16'h0580] = 8'h06;
    mem[16'h0581] = 8'h08;
    mem[16'h0582] = 8'h00;
    mem[16'h0583] = 8'h00;
    mem[16'h0584] = 8'h00;
    mem[16'h0585] = 8'h04; // PUSH RAX
    mem[16'h0586] = 8'h00;
    mem[16'h0587] = 8'h08; // POP RDI
    mem[16'h0588] = 8'h01;
    mem[16'h0589] = 8'h81; // ADDN RSP 8
    mem[16'h058A] = 8'h06;
    mem[16'h058B] = 8'h08;
    mem[16'h058C] = 8'h00;
    mem[16'h058D] = 8'h00;
    mem[16'h058E] = 8'h00;
    mem[16'h058F] = 8'h08; // POP RAX
    mem[16'h0590] = 8'h00;
    mem[16'h0591] = 8'h81; // ADDN RSP 8
    mem[16'h0592] = 8'h06;
    mem[16'h0593] = 8'h08;
    mem[16'h0594] = 8'h00;
    mem[16'h0595] = 8'h00;
    mem[16'h0596] = 8'h00;
    mem[16'h0597] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0598] = 8'h00;
    mem[16'h0599] = 8'h01;
    mem[16'h059A] = 8'h85; // SUBN RSP 8
    mem[16'h059B] = 8'h06;
    mem[16'h059C] = 8'h08;
    mem[16'h059D] = 8'h00;
    mem[16'h059E] = 8'h00;
    mem[16'h059F] = 8'h00;
    mem[16'h05A0] = 8'h04; // PUSH RDI
    mem[16'h05A1] = 8'h01;
    mem[16'h05A2] = 8'h81; // ADDN RSP 8
    mem[16'h05A3] = 8'h06;
    mem[16'h05A4] = 8'h08;
    mem[16'h05A5] = 8'h00;
    mem[16'h05A6] = 8'h00;
    mem[16'h05A7] = 8'h00;
    mem[16'h05A8] = 8'h22; // JMP .Lend3
    mem[16'h05A9] = 8'h01;
    mem[16'h05AA] = 8'h07;
    mem[16'h05AB] = 8'h00;
    mem[16'h05AC] = 8'h00;
    mem[16'h05AD] = 8'h00;
    mem[16'h05AE] = 8'h00;
    mem[16'h05AF] = 8'h00;
    mem[16'h05B0] = 8'h00;
                          // .Lelse3:
    mem[16'h05B1] = 8'h40; // MOV RAX RBP
    mem[16'h05B2] = 8'h00;
    mem[16'h05B3] = 8'h05;
    mem[16'h05B4] = 8'h85; // SUBN RAX 16
    mem[16'h05B5] = 8'h00;
    mem[16'h05B6] = 8'h10;
    mem[16'h05B7] = 8'h00;
    mem[16'h05B8] = 8'h00;
    mem[16'h05B9] = 8'h00;
    mem[16'h05BA] = 8'h85; // SUBN RSP 8
    mem[16'h05BB] = 8'h06;
    mem[16'h05BC] = 8'h08;
    mem[16'h05BD] = 8'h00;
    mem[16'h05BE] = 8'h00;
    mem[16'h05BF] = 8'h00;
    mem[16'h05C0] = 8'h04; // PUSH RAX
    mem[16'h05C1] = 8'h00;
    mem[16'h05C2] = 8'h85; // SUBN RSP 8
    mem[16'h05C3] = 8'h06;
    mem[16'h05C4] = 8'h08;
    mem[16'h05C5] = 8'h00;
    mem[16'h05C6] = 8'h00;
    mem[16'h05C7] = 8'h00;
    mem[16'h05C8] = 8'h05; // PUSHN 0
    mem[16'h05C9] = 8'h00;
    mem[16'h05CA] = 8'h00;
    mem[16'h05CB] = 8'h00;
    mem[16'h05CC] = 8'h00;
    mem[16'h05CD] = 8'h00;
    mem[16'h05CE] = 8'h08; // POP RDI
    mem[16'h05CF] = 8'h01;
    mem[16'h05D0] = 8'h81; // ADDN RSP 8
    mem[16'h05D1] = 8'h06;
    mem[16'h05D2] = 8'h08;
    mem[16'h05D3] = 8'h00;
    mem[16'h05D4] = 8'h00;
    mem[16'h05D5] = 8'h00;
    mem[16'h05D6] = 8'h08; // POP RAX
    mem[16'h05D7] = 8'h00;
    mem[16'h05D8] = 8'h81; // ADDN RSP 8
    mem[16'h05D9] = 8'h06;
    mem[16'h05DA] = 8'h08;
    mem[16'h05DB] = 8'h00;
    mem[16'h05DC] = 8'h00;
    mem[16'h05DD] = 8'h00;
    mem[16'h05DE] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h05DF] = 8'h00;
    mem[16'h05E0] = 8'h01;
    mem[16'h05E1] = 8'h85; // SUBN RSP 8
    mem[16'h05E2] = 8'h06;
    mem[16'h05E3] = 8'h08;
    mem[16'h05E4] = 8'h00;
    mem[16'h05E5] = 8'h00;
    mem[16'h05E6] = 8'h00;
    mem[16'h05E7] = 8'h04; // PUSH RDI
    mem[16'h05E8] = 8'h01;
    mem[16'h05E9] = 8'h81; // ADDN RSP 8
    mem[16'h05EA] = 8'h06;
    mem[16'h05EB] = 8'h08;
    mem[16'h05EC] = 8'h00;
    mem[16'h05ED] = 8'h00;
    mem[16'h05EE] = 8'h00;
    mem[16'h05EF] = 8'h40; // MOV RAX RBP
    mem[16'h05F0] = 8'h00;
    mem[16'h05F1] = 8'h05;
    mem[16'h05F2] = 8'h85; // SUBN RAX 12
    mem[16'h05F3] = 8'h00;
    mem[16'h05F4] = 8'h0C;
    mem[16'h05F5] = 8'h00;
    mem[16'h05F6] = 8'h00;
    mem[16'h05F7] = 8'h00;
    mem[16'h05F8] = 8'h85; // SUBN RSP 8
    mem[16'h05F9] = 8'h06;
    mem[16'h05FA] = 8'h08;
    mem[16'h05FB] = 8'h00;
    mem[16'h05FC] = 8'h00;
    mem[16'h05FD] = 8'h00;
    mem[16'h05FE] = 8'h04; // PUSH RAX
    mem[16'h05FF] = 8'h00;
    mem[16'h0600] = 8'h40; // MOV RAX RBP
    mem[16'h0601] = 8'h00;
    mem[16'h0602] = 8'h05;
    mem[16'h0603] = 8'h85; // SUBN RAX 28
    mem[16'h0604] = 8'h00;
    mem[16'h0605] = 8'h1C;
    mem[16'h0606] = 8'h00;
    mem[16'h0607] = 8'h00;
    mem[16'h0608] = 8'h00;
    mem[16'h0609] = 8'h85; // SUBN RSP 8
    mem[16'h060A] = 8'h06;
    mem[16'h060B] = 8'h08;
    mem[16'h060C] = 8'h00;
    mem[16'h060D] = 8'h00;
    mem[16'h060E] = 8'h00;
    mem[16'h060F] = 8'h04; // PUSH RAX
    mem[16'h0610] = 8'h00;
    mem[16'h0611] = 8'h08; // POP RAX
    mem[16'h0612] = 8'h00;
    mem[16'h0613] = 8'h81; // ADDN RSP 8
    mem[16'h0614] = 8'h06;
    mem[16'h0615] = 8'h08;
    mem[16'h0616] = 8'h00;
    mem[16'h0617] = 8'h00;
    mem[16'h0618] = 8'h00;
    mem[16'h0619] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h061A] = 8'h00;
    mem[16'h061B] = 8'h00;
    mem[16'h061C] = 8'h85; // SUBN RSP 8
    mem[16'h061D] = 8'h06;
    mem[16'h061E] = 8'h08;
    mem[16'h061F] = 8'h00;
    mem[16'h0620] = 8'h00;
    mem[16'h0621] = 8'h00;
    mem[16'h0622] = 8'h04; // PUSH RAX
    mem[16'h0623] = 8'h00;
    mem[16'h0624] = 8'h40; // MOV RAX RBP
    mem[16'h0625] = 8'h00;
    mem[16'h0626] = 8'h05;
    mem[16'h0627] = 8'h85; // SUBN RAX 32
    mem[16'h0628] = 8'h00;
    mem[16'h0629] = 8'h20;
    mem[16'h062A] = 8'h00;
    mem[16'h062B] = 8'h00;
    mem[16'h062C] = 8'h00;
    mem[16'h062D] = 8'h85; // SUBN RSP 8
    mem[16'h062E] = 8'h06;
    mem[16'h062F] = 8'h08;
    mem[16'h0630] = 8'h00;
    mem[16'h0631] = 8'h00;
    mem[16'h0632] = 8'h00;
    mem[16'h0633] = 8'h04; // PUSH RAX
    mem[16'h0634] = 8'h00;
    mem[16'h0635] = 8'h08; // POP RAX
    mem[16'h0636] = 8'h00;
    mem[16'h0637] = 8'h81; // ADDN RSP 8
    mem[16'h0638] = 8'h06;
    mem[16'h0639] = 8'h08;
    mem[16'h063A] = 8'h00;
    mem[16'h063B] = 8'h00;
    mem[16'h063C] = 8'h00;
    mem[16'h063D] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h063E] = 8'h00;
    mem[16'h063F] = 8'h00;
    mem[16'h0640] = 8'h85; // SUBN RSP 8
    mem[16'h0641] = 8'h06;
    mem[16'h0642] = 8'h08;
    mem[16'h0643] = 8'h00;
    mem[16'h0644] = 8'h00;
    mem[16'h0645] = 8'h00;
    mem[16'h0646] = 8'h04; // PUSH RAX
    mem[16'h0647] = 8'h00;
    mem[16'h0648] = 8'h08; // POP RDI
    mem[16'h0649] = 8'h01;
    mem[16'h064A] = 8'h81; // ADDN RSP 8
    mem[16'h064B] = 8'h06;
    mem[16'h064C] = 8'h08;
    mem[16'h064D] = 8'h00;
    mem[16'h064E] = 8'h00;
    mem[16'h064F] = 8'h00;
    mem[16'h0650] = 8'h08; // POP RAX
    mem[16'h0651] = 8'h00;
    mem[16'h0652] = 8'h81; // ADDN RSP 8
    mem[16'h0653] = 8'h06;
    mem[16'h0654] = 8'h08;
    mem[16'h0655] = 8'h00;
    mem[16'h0656] = 8'h00;
    mem[16'h0657] = 8'h00;
    mem[16'h0658] = 8'h84; // SUB RAX RDI
    mem[16'h0659] = 8'h00;
    mem[16'h065A] = 8'h01;
    mem[16'h065B] = 8'h85; // SUBN RSP 8
    mem[16'h065C] = 8'h06;
    mem[16'h065D] = 8'h08;
    mem[16'h065E] = 8'h00;
    mem[16'h065F] = 8'h00;
    mem[16'h0660] = 8'h00;
    mem[16'h0661] = 8'h04; // PUSH RAX
    mem[16'h0662] = 8'h00;
    mem[16'h0663] = 8'h08; // POP RDI
    mem[16'h0664] = 8'h01;
    mem[16'h0665] = 8'h81; // ADDN RSP 8
    mem[16'h0666] = 8'h06;
    mem[16'h0667] = 8'h08;
    mem[16'h0668] = 8'h00;
    mem[16'h0669] = 8'h00;
    mem[16'h066A] = 8'h00;
    mem[16'h066B] = 8'h08; // POP RAX
    mem[16'h066C] = 8'h00;
    mem[16'h066D] = 8'h81; // ADDN RSP 8
    mem[16'h066E] = 8'h06;
    mem[16'h066F] = 8'h08;
    mem[16'h0670] = 8'h00;
    mem[16'h0671] = 8'h00;
    mem[16'h0672] = 8'h00;
    mem[16'h0673] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0674] = 8'h00;
    mem[16'h0675] = 8'h01;
    mem[16'h0676] = 8'h85; // SUBN RSP 8
    mem[16'h0677] = 8'h06;
    mem[16'h0678] = 8'h08;
    mem[16'h0679] = 8'h00;
    mem[16'h067A] = 8'h00;
    mem[16'h067B] = 8'h00;
    mem[16'h067C] = 8'h04; // PUSH RDI
    mem[16'h067D] = 8'h01;
    mem[16'h067E] = 8'h81; // ADDN RSP 8
    mem[16'h067F] = 8'h06;
    mem[16'h0680] = 8'h08;
    mem[16'h0681] = 8'h00;
    mem[16'h0682] = 8'h00;
    mem[16'h0683] = 8'h00;
    mem[16'h0684] = 8'h40; // MOV RAX RBP
    mem[16'h0685] = 8'h00;
    mem[16'h0686] = 8'h05;
    mem[16'h0687] = 8'h85; // SUBN RAX 8
    mem[16'h0688] = 8'h00;
    mem[16'h0689] = 8'h08;
    mem[16'h068A] = 8'h00;
    mem[16'h068B] = 8'h00;
    mem[16'h068C] = 8'h00;
    mem[16'h068D] = 8'h85; // SUBN RSP 8
    mem[16'h068E] = 8'h06;
    mem[16'h068F] = 8'h08;
    mem[16'h0690] = 8'h00;
    mem[16'h0691] = 8'h00;
    mem[16'h0692] = 8'h00;
    mem[16'h0693] = 8'h04; // PUSH RAX
    mem[16'h0694] = 8'h00;
    mem[16'h0695] = 8'h85; // SUBN RSP 8
    mem[16'h0696] = 8'h06;
    mem[16'h0697] = 8'h08;
    mem[16'h0698] = 8'h00;
    mem[16'h0699] = 8'h00;
    mem[16'h069A] = 8'h00;
    mem[16'h069B] = 8'h05; // PUSHN 8
    mem[16'h069C] = 8'h00;
    mem[16'h069D] = 8'h08;
    mem[16'h069E] = 8'h00;
    mem[16'h069F] = 8'h00;
    mem[16'h06A0] = 8'h00;
    mem[16'h06A1] = 8'h40; // MOV RAX RBP
    mem[16'h06A2] = 8'h00;
    mem[16'h06A3] = 8'h05;
    mem[16'h06A4] = 8'h85; // SUBN RAX 12
    mem[16'h06A5] = 8'h00;
    mem[16'h06A6] = 8'h0C;
    mem[16'h06A7] = 8'h00;
    mem[16'h06A8] = 8'h00;
    mem[16'h06A9] = 8'h00;
    mem[16'h06AA] = 8'h85; // SUBN RSP 8
    mem[16'h06AB] = 8'h06;
    mem[16'h06AC] = 8'h08;
    mem[16'h06AD] = 8'h00;
    mem[16'h06AE] = 8'h00;
    mem[16'h06AF] = 8'h00;
    mem[16'h06B0] = 8'h04; // PUSH RAX
    mem[16'h06B1] = 8'h00;
    mem[16'h06B2] = 8'h08; // POP RAX
    mem[16'h06B3] = 8'h00;
    mem[16'h06B4] = 8'h81; // ADDN RSP 8
    mem[16'h06B5] = 8'h06;
    mem[16'h06B6] = 8'h08;
    mem[16'h06B7] = 8'h00;
    mem[16'h06B8] = 8'h00;
    mem[16'h06B9] = 8'h00;
    mem[16'h06BA] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h06BB] = 8'h00;
    mem[16'h06BC] = 8'h00;
    mem[16'h06BD] = 8'h85; // SUBN RSP 8
    mem[16'h06BE] = 8'h06;
    mem[16'h06BF] = 8'h08;
    mem[16'h06C0] = 8'h00;
    mem[16'h06C1] = 8'h00;
    mem[16'h06C2] = 8'h00;
    mem[16'h06C3] = 8'h04; // PUSH RAX
    mem[16'h06C4] = 8'h00;
    mem[16'h06C5] = 8'h08; // POP RDI
    mem[16'h06C6] = 8'h01;
    mem[16'h06C7] = 8'h81; // ADDN RSP 8
    mem[16'h06C8] = 8'h06;
    mem[16'h06C9] = 8'h08;
    mem[16'h06CA] = 8'h00;
    mem[16'h06CB] = 8'h00;
    mem[16'h06CC] = 8'h00;
    mem[16'h06CD] = 8'h08; // POP RAX
    mem[16'h06CE] = 8'h00;
    mem[16'h06CF] = 8'h81; // ADDN RSP 8
    mem[16'h06D0] = 8'h06;
    mem[16'h06D1] = 8'h08;
    mem[16'h06D2] = 8'h00;
    mem[16'h06D3] = 8'h00;
    mem[16'h06D4] = 8'h00;
    mem[16'h06D5] = 8'h84; // SUB RAX RDI
    mem[16'h06D6] = 8'h00;
    mem[16'h06D7] = 8'h01;
    mem[16'h06D8] = 8'h85; // SUBN RSP 8
    mem[16'h06D9] = 8'h06;
    mem[16'h06DA] = 8'h08;
    mem[16'h06DB] = 8'h00;
    mem[16'h06DC] = 8'h00;
    mem[16'h06DD] = 8'h00;
    mem[16'h06DE] = 8'h04; // PUSH RAX
    mem[16'h06DF] = 8'h00;
    mem[16'h06E0] = 8'h08; // POP RDI
    mem[16'h06E1] = 8'h01;
    mem[16'h06E2] = 8'h81; // ADDN RSP 8
    mem[16'h06E3] = 8'h06;
    mem[16'h06E4] = 8'h08;
    mem[16'h06E5] = 8'h00;
    mem[16'h06E6] = 8'h00;
    mem[16'h06E7] = 8'h00;
    mem[16'h06E8] = 8'h08; // POP RAX
    mem[16'h06E9] = 8'h00;
    mem[16'h06EA] = 8'h81; // ADDN RSP 8
    mem[16'h06EB] = 8'h06;
    mem[16'h06EC] = 8'h08;
    mem[16'h06ED] = 8'h00;
    mem[16'h06EE] = 8'h00;
    mem[16'h06EF] = 8'h00;
    mem[16'h06F0] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h06F1] = 8'h00;
    mem[16'h06F2] = 8'h01;
    mem[16'h06F3] = 8'h85; // SUBN RSP 8
    mem[16'h06F4] = 8'h06;
    mem[16'h06F5] = 8'h08;
    mem[16'h06F6] = 8'h00;
    mem[16'h06F7] = 8'h00;
    mem[16'h06F8] = 8'h00;
    mem[16'h06F9] = 8'h04; // PUSH RDI
    mem[16'h06FA] = 8'h01;
    mem[16'h06FB] = 8'h81; // ADDN RSP 8
    mem[16'h06FC] = 8'h06;
    mem[16'h06FD] = 8'h08;
    mem[16'h06FE] = 8'h00;
    mem[16'h06FF] = 8'h00;
    mem[16'h0700] = 8'h00;
                          // .Lend3:
    mem[16'h0701] = 8'h40; // MOV RAX RBP
    mem[16'h0702] = 8'h00;
    mem[16'h0703] = 8'h05;
    mem[16'h0704] = 8'h85; // SUBN RAX 4
    mem[16'h0705] = 8'h00;
    mem[16'h0706] = 8'h04;
    mem[16'h0707] = 8'h00;
    mem[16'h0708] = 8'h00;
    mem[16'h0709] = 8'h00;
    mem[16'h070A] = 8'h85; // SUBN RSP 8
    mem[16'h070B] = 8'h06;
    mem[16'h070C] = 8'h08;
    mem[16'h070D] = 8'h00;
    mem[16'h070E] = 8'h00;
    mem[16'h070F] = 8'h00;
    mem[16'h0710] = 8'h04; // PUSH RAX
    mem[16'h0711] = 8'h00;
    mem[16'h0712] = 8'h85; // SUBN RSP 8
    mem[16'h0713] = 8'h06;
    mem[16'h0714] = 8'h08;
    mem[16'h0715] = 8'h00;
    mem[16'h0716] = 8'h00;
    mem[16'h0717] = 8'h00;
    mem[16'h0718] = 8'h05; // PUSHN 0
    mem[16'h0719] = 8'h00;
    mem[16'h071A] = 8'h00;
    mem[16'h071B] = 8'h00;
    mem[16'h071C] = 8'h00;
    mem[16'h071D] = 8'h00;
    mem[16'h071E] = 8'h08; // POP RDI
    mem[16'h071F] = 8'h01;
    mem[16'h0720] = 8'h81; // ADDN RSP 8
    mem[16'h0721] = 8'h06;
    mem[16'h0722] = 8'h08;
    mem[16'h0723] = 8'h00;
    mem[16'h0724] = 8'h00;
    mem[16'h0725] = 8'h00;
    mem[16'h0726] = 8'h08; // POP RAX
    mem[16'h0727] = 8'h00;
    mem[16'h0728] = 8'h81; // ADDN RSP 8
    mem[16'h0729] = 8'h06;
    mem[16'h072A] = 8'h08;
    mem[16'h072B] = 8'h00;
    mem[16'h072C] = 8'h00;
    mem[16'h072D] = 8'h00;
    mem[16'h072E] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h072F] = 8'h00;
    mem[16'h0730] = 8'h01;
    mem[16'h0731] = 8'h85; // SUBN RSP 8
    mem[16'h0732] = 8'h06;
    mem[16'h0733] = 8'h08;
    mem[16'h0734] = 8'h00;
    mem[16'h0735] = 8'h00;
    mem[16'h0736] = 8'h00;
    mem[16'h0737] = 8'h04; // PUSH RDI
    mem[16'h0738] = 8'h01;
    mem[16'h0739] = 8'h81; // ADDN RSP 8
    mem[16'h073A] = 8'h06;
    mem[16'h073B] = 8'h08;
    mem[16'h073C] = 8'h00;
    mem[16'h073D] = 8'h00;
    mem[16'h073E] = 8'h00;
                          // .Lbegin4:
    mem[16'h073F] = 8'h40; // MOV RAX RBP
    mem[16'h0740] = 8'h00;
    mem[16'h0741] = 8'h05;
    mem[16'h0742] = 8'h85; // SUBN RAX 4
    mem[16'h0743] = 8'h00;
    mem[16'h0744] = 8'h04;
    mem[16'h0745] = 8'h00;
    mem[16'h0746] = 8'h00;
    mem[16'h0747] = 8'h00;
    mem[16'h0748] = 8'h85; // SUBN RSP 8
    mem[16'h0749] = 8'h06;
    mem[16'h074A] = 8'h08;
    mem[16'h074B] = 8'h00;
    mem[16'h074C] = 8'h00;
    mem[16'h074D] = 8'h00;
    mem[16'h074E] = 8'h04; // PUSH RAX
    mem[16'h074F] = 8'h00;
    mem[16'h0750] = 8'h08; // POP RAX
    mem[16'h0751] = 8'h00;
    mem[16'h0752] = 8'h81; // ADDN RSP 8
    mem[16'h0753] = 8'h06;
    mem[16'h0754] = 8'h08;
    mem[16'h0755] = 8'h00;
    mem[16'h0756] = 8'h00;
    mem[16'h0757] = 8'h00;
    mem[16'h0758] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0759] = 8'h00;
    mem[16'h075A] = 8'h00;
    mem[16'h075B] = 8'h85; // SUBN RSP 8
    mem[16'h075C] = 8'h06;
    mem[16'h075D] = 8'h08;
    mem[16'h075E] = 8'h00;
    mem[16'h075F] = 8'h00;
    mem[16'h0760] = 8'h00;
    mem[16'h0761] = 8'h04; // PUSH RAX
    mem[16'h0762] = 8'h00;
    mem[16'h0763] = 8'h40; // MOV RAX RBP
    mem[16'h0764] = 8'h00;
    mem[16'h0765] = 8'h05;
    mem[16'h0766] = 8'h85; // SUBN RAX 8
    mem[16'h0767] = 8'h00;
    mem[16'h0768] = 8'h08;
    mem[16'h0769] = 8'h00;
    mem[16'h076A] = 8'h00;
    mem[16'h076B] = 8'h00;
    mem[16'h076C] = 8'h85; // SUBN RSP 8
    mem[16'h076D] = 8'h06;
    mem[16'h076E] = 8'h08;
    mem[16'h076F] = 8'h00;
    mem[16'h0770] = 8'h00;
    mem[16'h0771] = 8'h00;
    mem[16'h0772] = 8'h04; // PUSH RAX
    mem[16'h0773] = 8'h00;
    mem[16'h0774] = 8'h08; // POP RAX
    mem[16'h0775] = 8'h00;
    mem[16'h0776] = 8'h81; // ADDN RSP 8
    mem[16'h0777] = 8'h06;
    mem[16'h0778] = 8'h08;
    mem[16'h0779] = 8'h00;
    mem[16'h077A] = 8'h00;
    mem[16'h077B] = 8'h00;
    mem[16'h077C] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h077D] = 8'h00;
    mem[16'h077E] = 8'h00;
    mem[16'h077F] = 8'h85; // SUBN RSP 8
    mem[16'h0780] = 8'h06;
    mem[16'h0781] = 8'h08;
    mem[16'h0782] = 8'h00;
    mem[16'h0783] = 8'h00;
    mem[16'h0784] = 8'h00;
    mem[16'h0785] = 8'h04; // PUSH RAX
    mem[16'h0786] = 8'h00;
    mem[16'h0787] = 8'h08; // POP RDI
    mem[16'h0788] = 8'h01;
    mem[16'h0789] = 8'h81; // ADDN RSP 8
    mem[16'h078A] = 8'h06;
    mem[16'h078B] = 8'h08;
    mem[16'h078C] = 8'h00;
    mem[16'h078D] = 8'h00;
    mem[16'h078E] = 8'h00;
    mem[16'h078F] = 8'h08; // POP RAX
    mem[16'h0790] = 8'h00;
    mem[16'h0791] = 8'h81; // ADDN RSP 8
    mem[16'h0792] = 8'h06;
    mem[16'h0793] = 8'h08;
    mem[16'h0794] = 8'h00;
    mem[16'h0795] = 8'h00;
    mem[16'h0796] = 8'h00;
    mem[16'h0797] = 8'h90; // CMP RAX RDI
    mem[16'h0798] = 8'h00;
    mem[16'h0799] = 8'h01;
    mem[16'h079A] = 8'h18; // SETL RAX
    mem[16'h079B] = 8'h00;
    mem[16'h079C] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h079D] = 8'h00;
    mem[16'h079E] = 8'h00;
    mem[16'h079F] = 8'h85; // SUBN RSP 8
    mem[16'h07A0] = 8'h06;
    mem[16'h07A1] = 8'h08;
    mem[16'h07A2] = 8'h00;
    mem[16'h07A3] = 8'h00;
    mem[16'h07A4] = 8'h00;
    mem[16'h07A5] = 8'h04; // PUSH RAX
    mem[16'h07A6] = 8'h00;
    mem[16'h07A7] = 8'h08; // POP RAX
    mem[16'h07A8] = 8'h00;
    mem[16'h07A9] = 8'h81; // ADDN RSP 8
    mem[16'h07AA] = 8'h06;
    mem[16'h07AB] = 8'h08;
    mem[16'h07AC] = 8'h00;
    mem[16'h07AD] = 8'h00;
    mem[16'h07AE] = 8'h00;
    mem[16'h07AF] = 8'h91; // CMPN RAX 0
    mem[16'h07B0] = 8'h00;
    mem[16'h07B1] = 8'h00;
    mem[16'h07B2] = 8'h00;
    mem[16'h07B3] = 8'h00;
    mem[16'h07B4] = 8'h00;
    mem[16'h07B5] = 8'h26; // JE .Lend4
    mem[16'h07B6] = 8'h7C;
    mem[16'h07B7] = 8'h0C;
    mem[16'h07B8] = 8'h00;
    mem[16'h07B9] = 8'h00;
    mem[16'h07BA] = 8'h00;
    mem[16'h07BB] = 8'h00;
    mem[16'h07BC] = 8'h00;
    mem[16'h07BD] = 8'h00;
    mem[16'h07BE] = 8'h40; // MOV RAX RBP
    mem[16'h07BF] = 8'h00;
    mem[16'h07C0] = 8'h05;
    mem[16'h07C1] = 8'h85; // SUBN RAX 20
    mem[16'h07C2] = 8'h00;
    mem[16'h07C3] = 8'h14;
    mem[16'h07C4] = 8'h00;
    mem[16'h07C5] = 8'h00;
    mem[16'h07C6] = 8'h00;
    mem[16'h07C7] = 8'h85; // SUBN RSP 8
    mem[16'h07C8] = 8'h06;
    mem[16'h07C9] = 8'h08;
    mem[16'h07CA] = 8'h00;
    mem[16'h07CB] = 8'h00;
    mem[16'h07CC] = 8'h00;
    mem[16'h07CD] = 8'h04; // PUSH RAX
    mem[16'h07CE] = 8'h00;
    mem[16'h07CF] = 8'h85; // SUBN RSP 8
    mem[16'h07D0] = 8'h06;
    mem[16'h07D1] = 8'h08;
    mem[16'h07D2] = 8'h00;
    mem[16'h07D3] = 8'h00;
    mem[16'h07D4] = 8'h00;
    mem[16'h07D5] = 8'h05; // PUSHN 0
    mem[16'h07D6] = 8'h00;
    mem[16'h07D7] = 8'h00;
    mem[16'h07D8] = 8'h00;
    mem[16'h07D9] = 8'h00;
    mem[16'h07DA] = 8'h00;
    mem[16'h07DB] = 8'h08; // POP RDI
    mem[16'h07DC] = 8'h01;
    mem[16'h07DD] = 8'h81; // ADDN RSP 8
    mem[16'h07DE] = 8'h06;
    mem[16'h07DF] = 8'h08;
    mem[16'h07E0] = 8'h00;
    mem[16'h07E1] = 8'h00;
    mem[16'h07E2] = 8'h00;
    mem[16'h07E3] = 8'h08; // POP RAX
    mem[16'h07E4] = 8'h00;
    mem[16'h07E5] = 8'h81; // ADDN RSP 8
    mem[16'h07E6] = 8'h06;
    mem[16'h07E7] = 8'h08;
    mem[16'h07E8] = 8'h00;
    mem[16'h07E9] = 8'h00;
    mem[16'h07EA] = 8'h00;
    mem[16'h07EB] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h07EC] = 8'h00;
    mem[16'h07ED] = 8'h01;
    mem[16'h07EE] = 8'h85; // SUBN RSP 8
    mem[16'h07EF] = 8'h06;
    mem[16'h07F0] = 8'h08;
    mem[16'h07F1] = 8'h00;
    mem[16'h07F2] = 8'h00;
    mem[16'h07F3] = 8'h00;
    mem[16'h07F4] = 8'h04; // PUSH RDI
    mem[16'h07F5] = 8'h01;
    mem[16'h07F6] = 8'h81; // ADDN RSP 8
    mem[16'h07F7] = 8'h06;
    mem[16'h07F8] = 8'h08;
    mem[16'h07F9] = 8'h00;
    mem[16'h07FA] = 8'h00;
    mem[16'h07FB] = 8'h00;
                          // .Lbegin5:
    mem[16'h07FC] = 8'h40; // MOV RAX RBP
    mem[16'h07FD] = 8'h00;
    mem[16'h07FE] = 8'h05;
    mem[16'h07FF] = 8'h85; // SUBN RAX 20
    mem[16'h0800] = 8'h00;
    mem[16'h0801] = 8'h14;
    mem[16'h0802] = 8'h00;
    mem[16'h0803] = 8'h00;
    mem[16'h0804] = 8'h00;
    mem[16'h0805] = 8'h85; // SUBN RSP 8
    mem[16'h0806] = 8'h06;
    mem[16'h0807] = 8'h08;
    mem[16'h0808] = 8'h00;
    mem[16'h0809] = 8'h00;
    mem[16'h080A] = 8'h00;
    mem[16'h080B] = 8'h04; // PUSH RAX
    mem[16'h080C] = 8'h00;
    mem[16'h080D] = 8'h08; // POP RAX
    mem[16'h080E] = 8'h00;
    mem[16'h080F] = 8'h81; // ADDN RSP 8
    mem[16'h0810] = 8'h06;
    mem[16'h0811] = 8'h08;
    mem[16'h0812] = 8'h00;
    mem[16'h0813] = 8'h00;
    mem[16'h0814] = 8'h00;
    mem[16'h0815] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0816] = 8'h00;
    mem[16'h0817] = 8'h00;
    mem[16'h0818] = 8'h85; // SUBN RSP 8
    mem[16'h0819] = 8'h06;
    mem[16'h081A] = 8'h08;
    mem[16'h081B] = 8'h00;
    mem[16'h081C] = 8'h00;
    mem[16'h081D] = 8'h00;
    mem[16'h081E] = 8'h04; // PUSH RAX
    mem[16'h081F] = 8'h00;
    mem[16'h0820] = 8'h40; // MOV RAX RBP
    mem[16'h0821] = 8'h00;
    mem[16'h0822] = 8'h05;
    mem[16'h0823] = 8'h85; // SUBN RAX 24
    mem[16'h0824] = 8'h00;
    mem[16'h0825] = 8'h18;
    mem[16'h0826] = 8'h00;
    mem[16'h0827] = 8'h00;
    mem[16'h0828] = 8'h00;
    mem[16'h0829] = 8'h85; // SUBN RSP 8
    mem[16'h082A] = 8'h06;
    mem[16'h082B] = 8'h08;
    mem[16'h082C] = 8'h00;
    mem[16'h082D] = 8'h00;
    mem[16'h082E] = 8'h00;
    mem[16'h082F] = 8'h04; // PUSH RAX
    mem[16'h0830] = 8'h00;
    mem[16'h0831] = 8'h08; // POP RAX
    mem[16'h0832] = 8'h00;
    mem[16'h0833] = 8'h81; // ADDN RSP 8
    mem[16'h0834] = 8'h06;
    mem[16'h0835] = 8'h08;
    mem[16'h0836] = 8'h00;
    mem[16'h0837] = 8'h00;
    mem[16'h0838] = 8'h00;
    mem[16'h0839] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h083A] = 8'h00;
    mem[16'h083B] = 8'h00;
    mem[16'h083C] = 8'h85; // SUBN RSP 8
    mem[16'h083D] = 8'h06;
    mem[16'h083E] = 8'h08;
    mem[16'h083F] = 8'h00;
    mem[16'h0840] = 8'h00;
    mem[16'h0841] = 8'h00;
    mem[16'h0842] = 8'h04; // PUSH RAX
    mem[16'h0843] = 8'h00;
    mem[16'h0844] = 8'h08; // POP RDI
    mem[16'h0845] = 8'h01;
    mem[16'h0846] = 8'h81; // ADDN RSP 8
    mem[16'h0847] = 8'h06;
    mem[16'h0848] = 8'h08;
    mem[16'h0849] = 8'h00;
    mem[16'h084A] = 8'h00;
    mem[16'h084B] = 8'h00;
    mem[16'h084C] = 8'h08; // POP RAX
    mem[16'h084D] = 8'h00;
    mem[16'h084E] = 8'h81; // ADDN RSP 8
    mem[16'h084F] = 8'h06;
    mem[16'h0850] = 8'h08;
    mem[16'h0851] = 8'h00;
    mem[16'h0852] = 8'h00;
    mem[16'h0853] = 8'h00;
    mem[16'h0854] = 8'h90; // CMP RAX RDI
    mem[16'h0855] = 8'h00;
    mem[16'h0856] = 8'h01;
    mem[16'h0857] = 8'h18; // SETL RAX
    mem[16'h0858] = 8'h00;
    mem[16'h0859] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h085A] = 8'h00;
    mem[16'h085B] = 8'h00;
    mem[16'h085C] = 8'h85; // SUBN RSP 8
    mem[16'h085D] = 8'h06;
    mem[16'h085E] = 8'h08;
    mem[16'h085F] = 8'h00;
    mem[16'h0860] = 8'h00;
    mem[16'h0861] = 8'h00;
    mem[16'h0862] = 8'h04; // PUSH RAX
    mem[16'h0863] = 8'h00;
    mem[16'h0864] = 8'h08; // POP RAX
    mem[16'h0865] = 8'h00;
    mem[16'h0866] = 8'h81; // ADDN RSP 8
    mem[16'h0867] = 8'h06;
    mem[16'h0868] = 8'h08;
    mem[16'h0869] = 8'h00;
    mem[16'h086A] = 8'h00;
    mem[16'h086B] = 8'h00;
    mem[16'h086C] = 8'h91; // CMPN RAX 0
    mem[16'h086D] = 8'h00;
    mem[16'h086E] = 8'h00;
    mem[16'h086F] = 8'h00;
    mem[16'h0870] = 8'h00;
    mem[16'h0871] = 8'h00;
    mem[16'h0872] = 8'h26; // JE .Lend5
    mem[16'h0873] = 8'hFC;
    mem[16'h0874] = 8'h0A;
    mem[16'h0875] = 8'h00;
    mem[16'h0876] = 8'h00;
    mem[16'h0877] = 8'h00;
    mem[16'h0878] = 8'h00;
    mem[16'h0879] = 8'h00;
    mem[16'h087A] = 8'h00;
    mem[16'h087B] = 8'h85; // SUBN RSP 8
    mem[16'h087C] = 8'h06;
    mem[16'h087D] = 8'h08;
    mem[16'h087E] = 8'h00;
    mem[16'h087F] = 8'h00;
    mem[16'h0880] = 8'h00;
    mem[16'h0881] = 8'h06; // PUSHA pos
    mem[16'h0882] = 8'h09;
    mem[16'h0883] = 8'h00;
    mem[16'h0884] = 8'h00;
    mem[16'h0885] = 8'h00;
    mem[16'h0886] = 8'h00;
    mem[16'h0887] = 8'h00;
    mem[16'h0888] = 8'h00;
    mem[16'h0889] = 8'h00;
    mem[16'h088A] = 8'h40; // MOV RAX RBP
    mem[16'h088B] = 8'h00;
    mem[16'h088C] = 8'h05;
    mem[16'h088D] = 8'h85; // SUBN RAX 20
    mem[16'h088E] = 8'h00;
    mem[16'h088F] = 8'h14;
    mem[16'h0890] = 8'h00;
    mem[16'h0891] = 8'h00;
    mem[16'h0892] = 8'h00;
    mem[16'h0893] = 8'h85; // SUBN RSP 8
    mem[16'h0894] = 8'h06;
    mem[16'h0895] = 8'h08;
    mem[16'h0896] = 8'h00;
    mem[16'h0897] = 8'h00;
    mem[16'h0898] = 8'h00;
    mem[16'h0899] = 8'h04; // PUSH RAX
    mem[16'h089A] = 8'h00;
    mem[16'h089B] = 8'h08; // POP RAX
    mem[16'h089C] = 8'h00;
    mem[16'h089D] = 8'h81; // ADDN RSP 8
    mem[16'h089E] = 8'h06;
    mem[16'h089F] = 8'h08;
    mem[16'h08A0] = 8'h00;
    mem[16'h08A1] = 8'h00;
    mem[16'h08A2] = 8'h00;
    mem[16'h08A3] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h08A4] = 8'h00;
    mem[16'h08A5] = 8'h00;
    mem[16'h08A6] = 8'h85; // SUBN RSP 8
    mem[16'h08A7] = 8'h06;
    mem[16'h08A8] = 8'h08;
    mem[16'h08A9] = 8'h00;
    mem[16'h08AA] = 8'h00;
    mem[16'h08AB] = 8'h00;
    mem[16'h08AC] = 8'h04; // PUSH RAX
    mem[16'h08AD] = 8'h00;
    mem[16'h08AE] = 8'h08; // POP RDI
    mem[16'h08AF] = 8'h01;
    mem[16'h08B0] = 8'h81; // ADDN RSP 8
    mem[16'h08B1] = 8'h06;
    mem[16'h08B2] = 8'h08;
    mem[16'h08B3] = 8'h00;
    mem[16'h08B4] = 8'h00;
    mem[16'h08B5] = 8'h00;
    mem[16'h08B6] = 8'h08; // POP RAX
    mem[16'h08B7] = 8'h00;
    mem[16'h08B8] = 8'h81; // ADDN RSP 8
    mem[16'h08B9] = 8'h06;
    mem[16'h08BA] = 8'h08;
    mem[16'h08BB] = 8'h00;
    mem[16'h08BC] = 8'h00;
    mem[16'h08BD] = 8'h00;
    mem[16'h08BE] = 8'h89; // MULN RDI 8
    mem[16'h08BF] = 8'h01;
    mem[16'h08C0] = 8'h08;
    mem[16'h08C1] = 8'h00;
    mem[16'h08C2] = 8'h00;
    mem[16'h08C3] = 8'h00;
    mem[16'h08C4] = 8'h80; // ADD RAX RDI
    mem[16'h08C5] = 8'h00;
    mem[16'h08C6] = 8'h01;
    mem[16'h08C7] = 8'h85; // SUBN RSP 8
    mem[16'h08C8] = 8'h06;
    mem[16'h08C9] = 8'h08;
    mem[16'h08CA] = 8'h00;
    mem[16'h08CB] = 8'h00;
    mem[16'h08CC] = 8'h00;
    mem[16'h08CD] = 8'h04; // PUSH RAX
    mem[16'h08CE] = 8'h00;
    mem[16'h08CF] = 8'h85; // SUBN RSP 8
    mem[16'h08D0] = 8'h06;
    mem[16'h08D1] = 8'h08;
    mem[16'h08D2] = 8'h00;
    mem[16'h08D3] = 8'h00;
    mem[16'h08D4] = 8'h00;
    mem[16'h08D5] = 8'h05; // PUSHN 0
    mem[16'h08D6] = 8'h00;
    mem[16'h08D7] = 8'h00;
    mem[16'h08D8] = 8'h00;
    mem[16'h08D9] = 8'h00;
    mem[16'h08DA] = 8'h00;
    mem[16'h08DB] = 8'h08; // POP RDI
    mem[16'h08DC] = 8'h01;
    mem[16'h08DD] = 8'h81; // ADDN RSP 8
    mem[16'h08DE] = 8'h06;
    mem[16'h08DF] = 8'h08;
    mem[16'h08E0] = 8'h00;
    mem[16'h08E1] = 8'h00;
    mem[16'h08E2] = 8'h00;
    mem[16'h08E3] = 8'h08; // POP RAX
    mem[16'h08E4] = 8'h00;
    mem[16'h08E5] = 8'h81; // ADDN RSP 8
    mem[16'h08E6] = 8'h06;
    mem[16'h08E7] = 8'h08;
    mem[16'h08E8] = 8'h00;
    mem[16'h08E9] = 8'h00;
    mem[16'h08EA] = 8'h00;
    mem[16'h08EB] = 8'h89; // MULN RDI 4
    mem[16'h08EC] = 8'h01;
    mem[16'h08ED] = 8'h04;
    mem[16'h08EE] = 8'h00;
    mem[16'h08EF] = 8'h00;
    mem[16'h08F0] = 8'h00;
    mem[16'h08F1] = 8'h80; // ADD RAX RDI
    mem[16'h08F2] = 8'h00;
    mem[16'h08F3] = 8'h01;
    mem[16'h08F4] = 8'h85; // SUBN RSP 8
    mem[16'h08F5] = 8'h06;
    mem[16'h08F6] = 8'h08;
    mem[16'h08F7] = 8'h00;
    mem[16'h08F8] = 8'h00;
    mem[16'h08F9] = 8'h00;
    mem[16'h08FA] = 8'h04; // PUSH RAX
    mem[16'h08FB] = 8'h00;
    mem[16'h08FC] = 8'h08; // POP RAX
    mem[16'h08FD] = 8'h00;
    mem[16'h08FE] = 8'h81; // ADDN RSP 8
    mem[16'h08FF] = 8'h06;
    mem[16'h0900] = 8'h08;
    mem[16'h0901] = 8'h00;
    mem[16'h0902] = 8'h00;
    mem[16'h0903] = 8'h00;
    mem[16'h0904] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0905] = 8'h00;
    mem[16'h0906] = 8'h00;
    mem[16'h0907] = 8'h85; // SUBN RSP 8
    mem[16'h0908] = 8'h06;
    mem[16'h0909] = 8'h08;
    mem[16'h090A] = 8'h00;
    mem[16'h090B] = 8'h00;
    mem[16'h090C] = 8'h00;
    mem[16'h090D] = 8'h04; // PUSH RAX
    mem[16'h090E] = 8'h00;
    mem[16'h090F] = 8'h40; // MOV RAX RBP
    mem[16'h0910] = 8'h00;
    mem[16'h0911] = 8'h05;
    mem[16'h0912] = 8'h85; // SUBN RAX 16
    mem[16'h0913] = 8'h00;
    mem[16'h0914] = 8'h10;
    mem[16'h0915] = 8'h00;
    mem[16'h0916] = 8'h00;
    mem[16'h0917] = 8'h00;
    mem[16'h0918] = 8'h85; // SUBN RSP 8
    mem[16'h0919] = 8'h06;
    mem[16'h091A] = 8'h08;
    mem[16'h091B] = 8'h00;
    mem[16'h091C] = 8'h00;
    mem[16'h091D] = 8'h00;
    mem[16'h091E] = 8'h04; // PUSH RAX
    mem[16'h091F] = 8'h00;
    mem[16'h0920] = 8'h08; // POP RAX
    mem[16'h0921] = 8'h00;
    mem[16'h0922] = 8'h81; // ADDN RSP 8
    mem[16'h0923] = 8'h06;
    mem[16'h0924] = 8'h08;
    mem[16'h0925] = 8'h00;
    mem[16'h0926] = 8'h00;
    mem[16'h0927] = 8'h00;
    mem[16'h0928] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0929] = 8'h00;
    mem[16'h092A] = 8'h00;
    mem[16'h092B] = 8'h85; // SUBN RSP 8
    mem[16'h092C] = 8'h06;
    mem[16'h092D] = 8'h08;
    mem[16'h092E] = 8'h00;
    mem[16'h092F] = 8'h00;
    mem[16'h0930] = 8'h00;
    mem[16'h0931] = 8'h04; // PUSH RAX
    mem[16'h0932] = 8'h00;
    mem[16'h0933] = 8'h08; // POP RDI
    mem[16'h0934] = 8'h01;
    mem[16'h0935] = 8'h81; // ADDN RSP 8
    mem[16'h0936] = 8'h06;
    mem[16'h0937] = 8'h08;
    mem[16'h0938] = 8'h00;
    mem[16'h0939] = 8'h00;
    mem[16'h093A] = 8'h00;
    mem[16'h093B] = 8'h08; // POP RAX
    mem[16'h093C] = 8'h00;
    mem[16'h093D] = 8'h81; // ADDN RSP 8
    mem[16'h093E] = 8'h06;
    mem[16'h093F] = 8'h08;
    mem[16'h0940] = 8'h00;
    mem[16'h0941] = 8'h00;
    mem[16'h0942] = 8'h00;
    mem[16'h0943] = 8'h90; // CMP RAX RDI
    mem[16'h0944] = 8'h00;
    mem[16'h0945] = 8'h01;
    mem[16'h0946] = 8'h10; // SETE RAX
    mem[16'h0947] = 8'h00;
    mem[16'h0948] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h0949] = 8'h00;
    mem[16'h094A] = 8'h00;
    mem[16'h094B] = 8'h85; // SUBN RSP 8
    mem[16'h094C] = 8'h06;
    mem[16'h094D] = 8'h08;
    mem[16'h094E] = 8'h00;
    mem[16'h094F] = 8'h00;
    mem[16'h0950] = 8'h00;
    mem[16'h0951] = 8'h04; // PUSH RAX
    mem[16'h0952] = 8'h00;
    mem[16'h0953] = 8'h08; // POP RAX
    mem[16'h0954] = 8'h00;
    mem[16'h0955] = 8'h81; // ADDN RSP 8
    mem[16'h0956] = 8'h06;
    mem[16'h0957] = 8'h08;
    mem[16'h0958] = 8'h00;
    mem[16'h0959] = 8'h00;
    mem[16'h095A] = 8'h00;
    mem[16'h095B] = 8'h91; // CMPN RAX 0
    mem[16'h095C] = 8'h00;
    mem[16'h095D] = 8'h00;
    mem[16'h095E] = 8'h00;
    mem[16'h095F] = 8'h00;
    mem[16'h0960] = 8'h00;
    mem[16'h0961] = 8'h26; // JE .Lend6
    mem[16'h0962] = 8'h76;
    mem[16'h0963] = 8'h0A;
    mem[16'h0964] = 8'h00;
    mem[16'h0965] = 8'h00;
    mem[16'h0966] = 8'h00;
    mem[16'h0967] = 8'h00;
    mem[16'h0968] = 8'h00;
    mem[16'h0969] = 8'h00;
    mem[16'h096A] = 8'h85; // SUBN RSP 8
    mem[16'h096B] = 8'h06;
    mem[16'h096C] = 8'h08;
    mem[16'h096D] = 8'h00;
    mem[16'h096E] = 8'h00;
    mem[16'h096F] = 8'h00;
    mem[16'h0970] = 8'h06; // PUSHA pos
    mem[16'h0971] = 8'h09;
    mem[16'h0972] = 8'h00;
    mem[16'h0973] = 8'h00;
    mem[16'h0974] = 8'h00;
    mem[16'h0975] = 8'h00;
    mem[16'h0976] = 8'h00;
    mem[16'h0977] = 8'h00;
    mem[16'h0978] = 8'h00;
    mem[16'h0979] = 8'h40; // MOV RAX RBP
    mem[16'h097A] = 8'h00;
    mem[16'h097B] = 8'h05;
    mem[16'h097C] = 8'h85; // SUBN RAX 20
    mem[16'h097D] = 8'h00;
    mem[16'h097E] = 8'h14;
    mem[16'h097F] = 8'h00;
    mem[16'h0980] = 8'h00;
    mem[16'h0981] = 8'h00;
    mem[16'h0982] = 8'h85; // SUBN RSP 8
    mem[16'h0983] = 8'h06;
    mem[16'h0984] = 8'h08;
    mem[16'h0985] = 8'h00;
    mem[16'h0986] = 8'h00;
    mem[16'h0987] = 8'h00;
    mem[16'h0988] = 8'h04; // PUSH RAX
    mem[16'h0989] = 8'h00;
    mem[16'h098A] = 8'h08; // POP RAX
    mem[16'h098B] = 8'h00;
    mem[16'h098C] = 8'h81; // ADDN RSP 8
    mem[16'h098D] = 8'h06;
    mem[16'h098E] = 8'h08;
    mem[16'h098F] = 8'h00;
    mem[16'h0990] = 8'h00;
    mem[16'h0991] = 8'h00;
    mem[16'h0992] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0993] = 8'h00;
    mem[16'h0994] = 8'h00;
    mem[16'h0995] = 8'h85; // SUBN RSP 8
    mem[16'h0996] = 8'h06;
    mem[16'h0997] = 8'h08;
    mem[16'h0998] = 8'h00;
    mem[16'h0999] = 8'h00;
    mem[16'h099A] = 8'h00;
    mem[16'h099B] = 8'h04; // PUSH RAX
    mem[16'h099C] = 8'h00;
    mem[16'h099D] = 8'h08; // POP RDI
    mem[16'h099E] = 8'h01;
    mem[16'h099F] = 8'h81; // ADDN RSP 8
    mem[16'h09A0] = 8'h06;
    mem[16'h09A1] = 8'h08;
    mem[16'h09A2] = 8'h00;
    mem[16'h09A3] = 8'h00;
    mem[16'h09A4] = 8'h00;
    mem[16'h09A5] = 8'h08; // POP RAX
    mem[16'h09A6] = 8'h00;
    mem[16'h09A7] = 8'h81; // ADDN RSP 8
    mem[16'h09A8] = 8'h06;
    mem[16'h09A9] = 8'h08;
    mem[16'h09AA] = 8'h00;
    mem[16'h09AB] = 8'h00;
    mem[16'h09AC] = 8'h00;
    mem[16'h09AD] = 8'h89; // MULN RDI 8
    mem[16'h09AE] = 8'h01;
    mem[16'h09AF] = 8'h08;
    mem[16'h09B0] = 8'h00;
    mem[16'h09B1] = 8'h00;
    mem[16'h09B2] = 8'h00;
    mem[16'h09B3] = 8'h80; // ADD RAX RDI
    mem[16'h09B4] = 8'h00;
    mem[16'h09B5] = 8'h01;
    mem[16'h09B6] = 8'h85; // SUBN RSP 8
    mem[16'h09B7] = 8'h06;
    mem[16'h09B8] = 8'h08;
    mem[16'h09B9] = 8'h00;
    mem[16'h09BA] = 8'h00;
    mem[16'h09BB] = 8'h00;
    mem[16'h09BC] = 8'h04; // PUSH RAX
    mem[16'h09BD] = 8'h00;
    mem[16'h09BE] = 8'h85; // SUBN RSP 8
    mem[16'h09BF] = 8'h06;
    mem[16'h09C0] = 8'h08;
    mem[16'h09C1] = 8'h00;
    mem[16'h09C2] = 8'h00;
    mem[16'h09C3] = 8'h00;
    mem[16'h09C4] = 8'h05; // PUSHN 1
    mem[16'h09C5] = 8'h00;
    mem[16'h09C6] = 8'h01;
    mem[16'h09C7] = 8'h00;
    mem[16'h09C8] = 8'h00;
    mem[16'h09C9] = 8'h00;
    mem[16'h09CA] = 8'h08; // POP RDI
    mem[16'h09CB] = 8'h01;
    mem[16'h09CC] = 8'h81; // ADDN RSP 8
    mem[16'h09CD] = 8'h06;
    mem[16'h09CE] = 8'h08;
    mem[16'h09CF] = 8'h00;
    mem[16'h09D0] = 8'h00;
    mem[16'h09D1] = 8'h00;
    mem[16'h09D2] = 8'h08; // POP RAX
    mem[16'h09D3] = 8'h00;
    mem[16'h09D4] = 8'h81; // ADDN RSP 8
    mem[16'h09D5] = 8'h06;
    mem[16'h09D6] = 8'h08;
    mem[16'h09D7] = 8'h00;
    mem[16'h09D8] = 8'h00;
    mem[16'h09D9] = 8'h00;
    mem[16'h09DA] = 8'h89; // MULN RDI 4
    mem[16'h09DB] = 8'h01;
    mem[16'h09DC] = 8'h04;
    mem[16'h09DD] = 8'h00;
    mem[16'h09DE] = 8'h00;
    mem[16'h09DF] = 8'h00;
    mem[16'h09E0] = 8'h80; // ADD RAX RDI
    mem[16'h09E1] = 8'h00;
    mem[16'h09E2] = 8'h01;
    mem[16'h09E3] = 8'h85; // SUBN RSP 8
    mem[16'h09E4] = 8'h06;
    mem[16'h09E5] = 8'h08;
    mem[16'h09E6] = 8'h00;
    mem[16'h09E7] = 8'h00;
    mem[16'h09E8] = 8'h00;
    mem[16'h09E9] = 8'h04; // PUSH RAX
    mem[16'h09EA] = 8'h00;
    mem[16'h09EB] = 8'h08; // POP RAX
    mem[16'h09EC] = 8'h00;
    mem[16'h09ED] = 8'h81; // ADDN RSP 8
    mem[16'h09EE] = 8'h06;
    mem[16'h09EF] = 8'h08;
    mem[16'h09F0] = 8'h00;
    mem[16'h09F1] = 8'h00;
    mem[16'h09F2] = 8'h00;
    mem[16'h09F3] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h09F4] = 8'h00;
    mem[16'h09F5] = 8'h00;
    mem[16'h09F6] = 8'h85; // SUBN RSP 8
    mem[16'h09F7] = 8'h06;
    mem[16'h09F8] = 8'h08;
    mem[16'h09F9] = 8'h00;
    mem[16'h09FA] = 8'h00;
    mem[16'h09FB] = 8'h00;
    mem[16'h09FC] = 8'h04; // PUSH RAX
    mem[16'h09FD] = 8'h00;
    mem[16'h09FE] = 8'h40; // MOV RAX RBP
    mem[16'h09FF] = 8'h00;
    mem[16'h0A00] = 8'h05;
    mem[16'h0A01] = 8'h85; // SUBN RAX 12
    mem[16'h0A02] = 8'h00;
    mem[16'h0A03] = 8'h0C;
    mem[16'h0A04] = 8'h00;
    mem[16'h0A05] = 8'h00;
    mem[16'h0A06] = 8'h00;
    mem[16'h0A07] = 8'h85; // SUBN RSP 8
    mem[16'h0A08] = 8'h06;
    mem[16'h0A09] = 8'h08;
    mem[16'h0A0A] = 8'h00;
    mem[16'h0A0B] = 8'h00;
    mem[16'h0A0C] = 8'h00;
    mem[16'h0A0D] = 8'h04; // PUSH RAX
    mem[16'h0A0E] = 8'h00;
    mem[16'h0A0F] = 8'h08; // POP RAX
    mem[16'h0A10] = 8'h00;
    mem[16'h0A11] = 8'h81; // ADDN RSP 8
    mem[16'h0A12] = 8'h06;
    mem[16'h0A13] = 8'h08;
    mem[16'h0A14] = 8'h00;
    mem[16'h0A15] = 8'h00;
    mem[16'h0A16] = 8'h00;
    mem[16'h0A17] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0A18] = 8'h00;
    mem[16'h0A19] = 8'h00;
    mem[16'h0A1A] = 8'h85; // SUBN RSP 8
    mem[16'h0A1B] = 8'h06;
    mem[16'h0A1C] = 8'h08;
    mem[16'h0A1D] = 8'h00;
    mem[16'h0A1E] = 8'h00;
    mem[16'h0A1F] = 8'h00;
    mem[16'h0A20] = 8'h04; // PUSH RAX
    mem[16'h0A21] = 8'h00;
    mem[16'h0A22] = 8'h08; // POP RDI
    mem[16'h0A23] = 8'h01;
    mem[16'h0A24] = 8'h81; // ADDN RSP 8
    mem[16'h0A25] = 8'h06;
    mem[16'h0A26] = 8'h08;
    mem[16'h0A27] = 8'h00;
    mem[16'h0A28] = 8'h00;
    mem[16'h0A29] = 8'h00;
    mem[16'h0A2A] = 8'h08; // POP RAX
    mem[16'h0A2B] = 8'h00;
    mem[16'h0A2C] = 8'h81; // ADDN RSP 8
    mem[16'h0A2D] = 8'h06;
    mem[16'h0A2E] = 8'h08;
    mem[16'h0A2F] = 8'h00;
    mem[16'h0A30] = 8'h00;
    mem[16'h0A31] = 8'h00;
    mem[16'h0A32] = 8'h90; // CMP RAX RDI
    mem[16'h0A33] = 8'h00;
    mem[16'h0A34] = 8'h01;
    mem[16'h0A35] = 8'h10; // SETE RAX
    mem[16'h0A36] = 8'h00;
    mem[16'h0A37] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h0A38] = 8'h00;
    mem[16'h0A39] = 8'h00;
    mem[16'h0A3A] = 8'h85; // SUBN RSP 8
    mem[16'h0A3B] = 8'h06;
    mem[16'h0A3C] = 8'h08;
    mem[16'h0A3D] = 8'h00;
    mem[16'h0A3E] = 8'h00;
    mem[16'h0A3F] = 8'h00;
    mem[16'h0A40] = 8'h04; // PUSH RAX
    mem[16'h0A41] = 8'h00;
    mem[16'h0A42] = 8'h08; // POP RAX
    mem[16'h0A43] = 8'h00;
    mem[16'h0A44] = 8'h81; // ADDN RSP 8
    mem[16'h0A45] = 8'h06;
    mem[16'h0A46] = 8'h08;
    mem[16'h0A47] = 8'h00;
    mem[16'h0A48] = 8'h00;
    mem[16'h0A49] = 8'h00;
    mem[16'h0A4A] = 8'h91; // CMPN RAX 0
    mem[16'h0A4B] = 8'h00;
    mem[16'h0A4C] = 8'h00;
    mem[16'h0A4D] = 8'h00;
    mem[16'h0A4E] = 8'h00;
    mem[16'h0A4F] = 8'h00;
    mem[16'h0A50] = 8'h26; // JE .Lend7
    mem[16'h0A51] = 8'h76;
    mem[16'h0A52] = 8'h0A;
    mem[16'h0A53] = 8'h00;
    mem[16'h0A54] = 8'h00;
    mem[16'h0A55] = 8'h00;
    mem[16'h0A56] = 8'h00;
    mem[16'h0A57] = 8'h00;
    mem[16'h0A58] = 8'h00;
    mem[16'h0A59] = 8'h85; // SUBN RSP 8
    mem[16'h0A5A] = 8'h06;
    mem[16'h0A5B] = 8'h08;
    mem[16'h0A5C] = 8'h00;
    mem[16'h0A5D] = 8'h00;
    mem[16'h0A5E] = 8'h00;
    mem[16'h0A5F] = 8'h05; // PUSHN 0
    mem[16'h0A60] = 8'h00;
    mem[16'h0A61] = 8'h00;
    mem[16'h0A62] = 8'h00;
    mem[16'h0A63] = 8'h00;
    mem[16'h0A64] = 8'h00;
    mem[16'h0A65] = 8'h08; // POP RAX
    mem[16'h0A66] = 8'h00;
    mem[16'h0A67] = 8'h81; // ADDN RSP 8
    mem[16'h0A68] = 8'h06;
    mem[16'h0A69] = 8'h08;
    mem[16'h0A6A] = 8'h00;
    mem[16'h0A6B] = 8'h00;
    mem[16'h0A6C] = 8'h00;
    mem[16'h0A6D] = 8'h22; // JMP .Lreturn.check
    mem[16'h0A6E] = 8'h08;
    mem[16'h0A6F] = 8'h16;
    mem[16'h0A70] = 8'h00;
    mem[16'h0A71] = 8'h00;
    mem[16'h0A72] = 8'h00;
    mem[16'h0A73] = 8'h00;
    mem[16'h0A74] = 8'h00;
    mem[16'h0A75] = 8'h00;
                          // .Lend7:
                          // .Lend6:
    mem[16'h0A76] = 8'h40; // MOV RAX RBP
    mem[16'h0A77] = 8'h00;
    mem[16'h0A78] = 8'h05;
    mem[16'h0A79] = 8'h85; // SUBN RAX 20
    mem[16'h0A7A] = 8'h00;
    mem[16'h0A7B] = 8'h14;
    mem[16'h0A7C] = 8'h00;
    mem[16'h0A7D] = 8'h00;
    mem[16'h0A7E] = 8'h00;
    mem[16'h0A7F] = 8'h85; // SUBN RSP 8
    mem[16'h0A80] = 8'h06;
    mem[16'h0A81] = 8'h08;
    mem[16'h0A82] = 8'h00;
    mem[16'h0A83] = 8'h00;
    mem[16'h0A84] = 8'h00;
    mem[16'h0A85] = 8'h04; // PUSH RAX
    mem[16'h0A86] = 8'h00;
    mem[16'h0A87] = 8'h40; // MOV RAX RBP
    mem[16'h0A88] = 8'h00;
    mem[16'h0A89] = 8'h05;
    mem[16'h0A8A] = 8'h85; // SUBN RAX 20
    mem[16'h0A8B] = 8'h00;
    mem[16'h0A8C] = 8'h14;
    mem[16'h0A8D] = 8'h00;
    mem[16'h0A8E] = 8'h00;
    mem[16'h0A8F] = 8'h00;
    mem[16'h0A90] = 8'h85; // SUBN RSP 8
    mem[16'h0A91] = 8'h06;
    mem[16'h0A92] = 8'h08;
    mem[16'h0A93] = 8'h00;
    mem[16'h0A94] = 8'h00;
    mem[16'h0A95] = 8'h00;
    mem[16'h0A96] = 8'h04; // PUSH RAX
    mem[16'h0A97] = 8'h00;
    mem[16'h0A98] = 8'h08; // POP RAX
    mem[16'h0A99] = 8'h00;
    mem[16'h0A9A] = 8'h81; // ADDN RSP 8
    mem[16'h0A9B] = 8'h06;
    mem[16'h0A9C] = 8'h08;
    mem[16'h0A9D] = 8'h00;
    mem[16'h0A9E] = 8'h00;
    mem[16'h0A9F] = 8'h00;
    mem[16'h0AA0] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0AA1] = 8'h00;
    mem[16'h0AA2] = 8'h00;
    mem[16'h0AA3] = 8'h85; // SUBN RSP 8
    mem[16'h0AA4] = 8'h06;
    mem[16'h0AA5] = 8'h08;
    mem[16'h0AA6] = 8'h00;
    mem[16'h0AA7] = 8'h00;
    mem[16'h0AA8] = 8'h00;
    mem[16'h0AA9] = 8'h04; // PUSH RAX
    mem[16'h0AAA] = 8'h00;
    mem[16'h0AAB] = 8'h85; // SUBN RSP 8
    mem[16'h0AAC] = 8'h06;
    mem[16'h0AAD] = 8'h08;
    mem[16'h0AAE] = 8'h00;
    mem[16'h0AAF] = 8'h00;
    mem[16'h0AB0] = 8'h00;
    mem[16'h0AB1] = 8'h05; // PUSHN 1
    mem[16'h0AB2] = 8'h00;
    mem[16'h0AB3] = 8'h01;
    mem[16'h0AB4] = 8'h00;
    mem[16'h0AB5] = 8'h00;
    mem[16'h0AB6] = 8'h00;
    mem[16'h0AB7] = 8'h08; // POP RDI
    mem[16'h0AB8] = 8'h01;
    mem[16'h0AB9] = 8'h81; // ADDN RSP 8
    mem[16'h0ABA] = 8'h06;
    mem[16'h0ABB] = 8'h08;
    mem[16'h0ABC] = 8'h00;
    mem[16'h0ABD] = 8'h00;
    mem[16'h0ABE] = 8'h00;
    mem[16'h0ABF] = 8'h08; // POP RAX
    mem[16'h0AC0] = 8'h00;
    mem[16'h0AC1] = 8'h81; // ADDN RSP 8
    mem[16'h0AC2] = 8'h06;
    mem[16'h0AC3] = 8'h08;
    mem[16'h0AC4] = 8'h00;
    mem[16'h0AC5] = 8'h00;
    mem[16'h0AC6] = 8'h00;
    mem[16'h0AC7] = 8'h80; // ADD RAX RDI
    mem[16'h0AC8] = 8'h00;
    mem[16'h0AC9] = 8'h01;
    mem[16'h0ACA] = 8'h85; // SUBN RSP 8
    mem[16'h0ACB] = 8'h06;
    mem[16'h0ACC] = 8'h08;
    mem[16'h0ACD] = 8'h00;
    mem[16'h0ACE] = 8'h00;
    mem[16'h0ACF] = 8'h00;
    mem[16'h0AD0] = 8'h04; // PUSH RAX
    mem[16'h0AD1] = 8'h00;
    mem[16'h0AD2] = 8'h08; // POP RDI
    mem[16'h0AD3] = 8'h01;
    mem[16'h0AD4] = 8'h81; // ADDN RSP 8
    mem[16'h0AD5] = 8'h06;
    mem[16'h0AD6] = 8'h08;
    mem[16'h0AD7] = 8'h00;
    mem[16'h0AD8] = 8'h00;
    mem[16'h0AD9] = 8'h00;
    mem[16'h0ADA] = 8'h08; // POP RAX
    mem[16'h0ADB] = 8'h00;
    mem[16'h0ADC] = 8'h81; // ADDN RSP 8
    mem[16'h0ADD] = 8'h06;
    mem[16'h0ADE] = 8'h08;
    mem[16'h0ADF] = 8'h00;
    mem[16'h0AE0] = 8'h00;
    mem[16'h0AE1] = 8'h00;
    mem[16'h0AE2] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0AE3] = 8'h00;
    mem[16'h0AE4] = 8'h01;
    mem[16'h0AE5] = 8'h85; // SUBN RSP 8
    mem[16'h0AE6] = 8'h06;
    mem[16'h0AE7] = 8'h08;
    mem[16'h0AE8] = 8'h00;
    mem[16'h0AE9] = 8'h00;
    mem[16'h0AEA] = 8'h00;
    mem[16'h0AEB] = 8'h04; // PUSH RDI
    mem[16'h0AEC] = 8'h01;
    mem[16'h0AED] = 8'h81; // ADDN RSP 8
    mem[16'h0AEE] = 8'h06;
    mem[16'h0AEF] = 8'h08;
    mem[16'h0AF0] = 8'h00;
    mem[16'h0AF1] = 8'h00;
    mem[16'h0AF2] = 8'h00;
    mem[16'h0AF3] = 8'h22; // JMP .Lbegin5
    mem[16'h0AF4] = 8'hFC;
    mem[16'h0AF5] = 8'h07;
    mem[16'h0AF6] = 8'h00;
    mem[16'h0AF7] = 8'h00;
    mem[16'h0AF8] = 8'h00;
    mem[16'h0AF9] = 8'h00;
    mem[16'h0AFA] = 8'h00;
    mem[16'h0AFB] = 8'h00;
                          // .Lend5:
    mem[16'h0AFC] = 8'h40; // MOV RAX RBP
    mem[16'h0AFD] = 8'h00;
    mem[16'h0AFE] = 8'h05;
    mem[16'h0AFF] = 8'h85; // SUBN RAX 16
    mem[16'h0B00] = 8'h00;
    mem[16'h0B01] = 8'h10;
    mem[16'h0B02] = 8'h00;
    mem[16'h0B03] = 8'h00;
    mem[16'h0B04] = 8'h00;
    mem[16'h0B05] = 8'h85; // SUBN RSP 8
    mem[16'h0B06] = 8'h06;
    mem[16'h0B07] = 8'h08;
    mem[16'h0B08] = 8'h00;
    mem[16'h0B09] = 8'h00;
    mem[16'h0B0A] = 8'h00;
    mem[16'h0B0B] = 8'h04; // PUSH RAX
    mem[16'h0B0C] = 8'h00;
    mem[16'h0B0D] = 8'h40; // MOV RAX RBP
    mem[16'h0B0E] = 8'h00;
    mem[16'h0B0F] = 8'h05;
    mem[16'h0B10] = 8'h85; // SUBN RAX 16
    mem[16'h0B11] = 8'h00;
    mem[16'h0B12] = 8'h10;
    mem[16'h0B13] = 8'h00;
    mem[16'h0B14] = 8'h00;
    mem[16'h0B15] = 8'h00;
    mem[16'h0B16] = 8'h85; // SUBN RSP 8
    mem[16'h0B17] = 8'h06;
    mem[16'h0B18] = 8'h08;
    mem[16'h0B19] = 8'h00;
    mem[16'h0B1A] = 8'h00;
    mem[16'h0B1B] = 8'h00;
    mem[16'h0B1C] = 8'h04; // PUSH RAX
    mem[16'h0B1D] = 8'h00;
    mem[16'h0B1E] = 8'h08; // POP RAX
    mem[16'h0B1F] = 8'h00;
    mem[16'h0B20] = 8'h81; // ADDN RSP 8
    mem[16'h0B21] = 8'h06;
    mem[16'h0B22] = 8'h08;
    mem[16'h0B23] = 8'h00;
    mem[16'h0B24] = 8'h00;
    mem[16'h0B25] = 8'h00;
    mem[16'h0B26] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0B27] = 8'h00;
    mem[16'h0B28] = 8'h00;
    mem[16'h0B29] = 8'h85; // SUBN RSP 8
    mem[16'h0B2A] = 8'h06;
    mem[16'h0B2B] = 8'h08;
    mem[16'h0B2C] = 8'h00;
    mem[16'h0B2D] = 8'h00;
    mem[16'h0B2E] = 8'h00;
    mem[16'h0B2F] = 8'h04; // PUSH RAX
    mem[16'h0B30] = 8'h00;
    mem[16'h0B31] = 8'h85; // SUBN RSP 8
    mem[16'h0B32] = 8'h06;
    mem[16'h0B33] = 8'h08;
    mem[16'h0B34] = 8'h00;
    mem[16'h0B35] = 8'h00;
    mem[16'h0B36] = 8'h00;
    mem[16'h0B37] = 8'h05; // PUSHN 1
    mem[16'h0B38] = 8'h00;
    mem[16'h0B39] = 8'h01;
    mem[16'h0B3A] = 8'h00;
    mem[16'h0B3B] = 8'h00;
    mem[16'h0B3C] = 8'h00;
    mem[16'h0B3D] = 8'h08; // POP RDI
    mem[16'h0B3E] = 8'h01;
    mem[16'h0B3F] = 8'h81; // ADDN RSP 8
    mem[16'h0B40] = 8'h06;
    mem[16'h0B41] = 8'h08;
    mem[16'h0B42] = 8'h00;
    mem[16'h0B43] = 8'h00;
    mem[16'h0B44] = 8'h00;
    mem[16'h0B45] = 8'h08; // POP RAX
    mem[16'h0B46] = 8'h00;
    mem[16'h0B47] = 8'h81; // ADDN RSP 8
    mem[16'h0B48] = 8'h06;
    mem[16'h0B49] = 8'h08;
    mem[16'h0B4A] = 8'h00;
    mem[16'h0B4B] = 8'h00;
    mem[16'h0B4C] = 8'h00;
    mem[16'h0B4D] = 8'h80; // ADD RAX RDI
    mem[16'h0B4E] = 8'h00;
    mem[16'h0B4F] = 8'h01;
    mem[16'h0B50] = 8'h85; // SUBN RSP 8
    mem[16'h0B51] = 8'h06;
    mem[16'h0B52] = 8'h08;
    mem[16'h0B53] = 8'h00;
    mem[16'h0B54] = 8'h00;
    mem[16'h0B55] = 8'h00;
    mem[16'h0B56] = 8'h04; // PUSH RAX
    mem[16'h0B57] = 8'h00;
    mem[16'h0B58] = 8'h08; // POP RDI
    mem[16'h0B59] = 8'h01;
    mem[16'h0B5A] = 8'h81; // ADDN RSP 8
    mem[16'h0B5B] = 8'h06;
    mem[16'h0B5C] = 8'h08;
    mem[16'h0B5D] = 8'h00;
    mem[16'h0B5E] = 8'h00;
    mem[16'h0B5F] = 8'h00;
    mem[16'h0B60] = 8'h08; // POP RAX
    mem[16'h0B61] = 8'h00;
    mem[16'h0B62] = 8'h81; // ADDN RSP 8
    mem[16'h0B63] = 8'h06;
    mem[16'h0B64] = 8'h08;
    mem[16'h0B65] = 8'h00;
    mem[16'h0B66] = 8'h00;
    mem[16'h0B67] = 8'h00;
    mem[16'h0B68] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0B69] = 8'h00;
    mem[16'h0B6A] = 8'h01;
    mem[16'h0B6B] = 8'h85; // SUBN RSP 8
    mem[16'h0B6C] = 8'h06;
    mem[16'h0B6D] = 8'h08;
    mem[16'h0B6E] = 8'h00;
    mem[16'h0B6F] = 8'h00;
    mem[16'h0B70] = 8'h00;
    mem[16'h0B71] = 8'h04; // PUSH RDI
    mem[16'h0B72] = 8'h01;
    mem[16'h0B73] = 8'h81; // ADDN RSP 8
    mem[16'h0B74] = 8'h06;
    mem[16'h0B75] = 8'h08;
    mem[16'h0B76] = 8'h00;
    mem[16'h0B77] = 8'h00;
    mem[16'h0B78] = 8'h00;
    mem[16'h0B79] = 8'h40; // MOV RAX RBP
    mem[16'h0B7A] = 8'h00;
    mem[16'h0B7B] = 8'h05;
    mem[16'h0B7C] = 8'h85; // SUBN RAX 12
    mem[16'h0B7D] = 8'h00;
    mem[16'h0B7E] = 8'h0C;
    mem[16'h0B7F] = 8'h00;
    mem[16'h0B80] = 8'h00;
    mem[16'h0B81] = 8'h00;
    mem[16'h0B82] = 8'h85; // SUBN RSP 8
    mem[16'h0B83] = 8'h06;
    mem[16'h0B84] = 8'h08;
    mem[16'h0B85] = 8'h00;
    mem[16'h0B86] = 8'h00;
    mem[16'h0B87] = 8'h00;
    mem[16'h0B88] = 8'h04; // PUSH RAX
    mem[16'h0B89] = 8'h00;
    mem[16'h0B8A] = 8'h40; // MOV RAX RBP
    mem[16'h0B8B] = 8'h00;
    mem[16'h0B8C] = 8'h05;
    mem[16'h0B8D] = 8'h85; // SUBN RAX 12
    mem[16'h0B8E] = 8'h00;
    mem[16'h0B8F] = 8'h0C;
    mem[16'h0B90] = 8'h00;
    mem[16'h0B91] = 8'h00;
    mem[16'h0B92] = 8'h00;
    mem[16'h0B93] = 8'h85; // SUBN RSP 8
    mem[16'h0B94] = 8'h06;
    mem[16'h0B95] = 8'h08;
    mem[16'h0B96] = 8'h00;
    mem[16'h0B97] = 8'h00;
    mem[16'h0B98] = 8'h00;
    mem[16'h0B99] = 8'h04; // PUSH RAX
    mem[16'h0B9A] = 8'h00;
    mem[16'h0B9B] = 8'h08; // POP RAX
    mem[16'h0B9C] = 8'h00;
    mem[16'h0B9D] = 8'h81; // ADDN RSP 8
    mem[16'h0B9E] = 8'h06;
    mem[16'h0B9F] = 8'h08;
    mem[16'h0BA0] = 8'h00;
    mem[16'h0BA1] = 8'h00;
    mem[16'h0BA2] = 8'h00;
    mem[16'h0BA3] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0BA4] = 8'h00;
    mem[16'h0BA5] = 8'h00;
    mem[16'h0BA6] = 8'h85; // SUBN RSP 8
    mem[16'h0BA7] = 8'h06;
    mem[16'h0BA8] = 8'h08;
    mem[16'h0BA9] = 8'h00;
    mem[16'h0BAA] = 8'h00;
    mem[16'h0BAB] = 8'h00;
    mem[16'h0BAC] = 8'h04; // PUSH RAX
    mem[16'h0BAD] = 8'h00;
    mem[16'h0BAE] = 8'h85; // SUBN RSP 8
    mem[16'h0BAF] = 8'h06;
    mem[16'h0BB0] = 8'h08;
    mem[16'h0BB1] = 8'h00;
    mem[16'h0BB2] = 8'h00;
    mem[16'h0BB3] = 8'h00;
    mem[16'h0BB4] = 8'h05; // PUSHN 1
    mem[16'h0BB5] = 8'h00;
    mem[16'h0BB6] = 8'h01;
    mem[16'h0BB7] = 8'h00;
    mem[16'h0BB8] = 8'h00;
    mem[16'h0BB9] = 8'h00;
    mem[16'h0BBA] = 8'h08; // POP RDI
    mem[16'h0BBB] = 8'h01;
    mem[16'h0BBC] = 8'h81; // ADDN RSP 8
    mem[16'h0BBD] = 8'h06;
    mem[16'h0BBE] = 8'h08;
    mem[16'h0BBF] = 8'h00;
    mem[16'h0BC0] = 8'h00;
    mem[16'h0BC1] = 8'h00;
    mem[16'h0BC2] = 8'h08; // POP RAX
    mem[16'h0BC3] = 8'h00;
    mem[16'h0BC4] = 8'h81; // ADDN RSP 8
    mem[16'h0BC5] = 8'h06;
    mem[16'h0BC6] = 8'h08;
    mem[16'h0BC7] = 8'h00;
    mem[16'h0BC8] = 8'h00;
    mem[16'h0BC9] = 8'h00;
    mem[16'h0BCA] = 8'h80; // ADD RAX RDI
    mem[16'h0BCB] = 8'h00;
    mem[16'h0BCC] = 8'h01;
    mem[16'h0BCD] = 8'h85; // SUBN RSP 8
    mem[16'h0BCE] = 8'h06;
    mem[16'h0BCF] = 8'h08;
    mem[16'h0BD0] = 8'h00;
    mem[16'h0BD1] = 8'h00;
    mem[16'h0BD2] = 8'h00;
    mem[16'h0BD3] = 8'h04; // PUSH RAX
    mem[16'h0BD4] = 8'h00;
    mem[16'h0BD5] = 8'h08; // POP RDI
    mem[16'h0BD6] = 8'h01;
    mem[16'h0BD7] = 8'h81; // ADDN RSP 8
    mem[16'h0BD8] = 8'h06;
    mem[16'h0BD9] = 8'h08;
    mem[16'h0BDA] = 8'h00;
    mem[16'h0BDB] = 8'h00;
    mem[16'h0BDC] = 8'h00;
    mem[16'h0BDD] = 8'h08; // POP RAX
    mem[16'h0BDE] = 8'h00;
    mem[16'h0BDF] = 8'h81; // ADDN RSP 8
    mem[16'h0BE0] = 8'h06;
    mem[16'h0BE1] = 8'h08;
    mem[16'h0BE2] = 8'h00;
    mem[16'h0BE3] = 8'h00;
    mem[16'h0BE4] = 8'h00;
    mem[16'h0BE5] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0BE6] = 8'h00;
    mem[16'h0BE7] = 8'h01;
    mem[16'h0BE8] = 8'h85; // SUBN RSP 8
    mem[16'h0BE9] = 8'h06;
    mem[16'h0BEA] = 8'h08;
    mem[16'h0BEB] = 8'h00;
    mem[16'h0BEC] = 8'h00;
    mem[16'h0BED] = 8'h00;
    mem[16'h0BEE] = 8'h04; // PUSH RDI
    mem[16'h0BEF] = 8'h01;
    mem[16'h0BF0] = 8'h81; // ADDN RSP 8
    mem[16'h0BF1] = 8'h06;
    mem[16'h0BF2] = 8'h08;
    mem[16'h0BF3] = 8'h00;
    mem[16'h0BF4] = 8'h00;
    mem[16'h0BF5] = 8'h00;
    mem[16'h0BF6] = 8'h40; // MOV RAX RBP
    mem[16'h0BF7] = 8'h00;
    mem[16'h0BF8] = 8'h05;
    mem[16'h0BF9] = 8'h85; // SUBN RAX 4
    mem[16'h0BFA] = 8'h00;
    mem[16'h0BFB] = 8'h04;
    mem[16'h0BFC] = 8'h00;
    mem[16'h0BFD] = 8'h00;
    mem[16'h0BFE] = 8'h00;
    mem[16'h0BFF] = 8'h85; // SUBN RSP 8
    mem[16'h0C00] = 8'h06;
    mem[16'h0C01] = 8'h08;
    mem[16'h0C02] = 8'h00;
    mem[16'h0C03] = 8'h00;
    mem[16'h0C04] = 8'h00;
    mem[16'h0C05] = 8'h04; // PUSH RAX
    mem[16'h0C06] = 8'h00;
    mem[16'h0C07] = 8'h40; // MOV RAX RBP
    mem[16'h0C08] = 8'h00;
    mem[16'h0C09] = 8'h05;
    mem[16'h0C0A] = 8'h85; // SUBN RAX 4
    mem[16'h0C0B] = 8'h00;
    mem[16'h0C0C] = 8'h04;
    mem[16'h0C0D] = 8'h00;
    mem[16'h0C0E] = 8'h00;
    mem[16'h0C0F] = 8'h00;
    mem[16'h0C10] = 8'h85; // SUBN RSP 8
    mem[16'h0C11] = 8'h06;
    mem[16'h0C12] = 8'h08;
    mem[16'h0C13] = 8'h00;
    mem[16'h0C14] = 8'h00;
    mem[16'h0C15] = 8'h00;
    mem[16'h0C16] = 8'h04; // PUSH RAX
    mem[16'h0C17] = 8'h00;
    mem[16'h0C18] = 8'h08; // POP RAX
    mem[16'h0C19] = 8'h00;
    mem[16'h0C1A] = 8'h81; // ADDN RSP 8
    mem[16'h0C1B] = 8'h06;
    mem[16'h0C1C] = 8'h08;
    mem[16'h0C1D] = 8'h00;
    mem[16'h0C1E] = 8'h00;
    mem[16'h0C1F] = 8'h00;
    mem[16'h0C20] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0C21] = 8'h00;
    mem[16'h0C22] = 8'h00;
    mem[16'h0C23] = 8'h85; // SUBN RSP 8
    mem[16'h0C24] = 8'h06;
    mem[16'h0C25] = 8'h08;
    mem[16'h0C26] = 8'h00;
    mem[16'h0C27] = 8'h00;
    mem[16'h0C28] = 8'h00;
    mem[16'h0C29] = 8'h04; // PUSH RAX
    mem[16'h0C2A] = 8'h00;
    mem[16'h0C2B] = 8'h85; // SUBN RSP 8
    mem[16'h0C2C] = 8'h06;
    mem[16'h0C2D] = 8'h08;
    mem[16'h0C2E] = 8'h00;
    mem[16'h0C2F] = 8'h00;
    mem[16'h0C30] = 8'h00;
    mem[16'h0C31] = 8'h05; // PUSHN 1
    mem[16'h0C32] = 8'h00;
    mem[16'h0C33] = 8'h01;
    mem[16'h0C34] = 8'h00;
    mem[16'h0C35] = 8'h00;
    mem[16'h0C36] = 8'h00;
    mem[16'h0C37] = 8'h08; // POP RDI
    mem[16'h0C38] = 8'h01;
    mem[16'h0C39] = 8'h81; // ADDN RSP 8
    mem[16'h0C3A] = 8'h06;
    mem[16'h0C3B] = 8'h08;
    mem[16'h0C3C] = 8'h00;
    mem[16'h0C3D] = 8'h00;
    mem[16'h0C3E] = 8'h00;
    mem[16'h0C3F] = 8'h08; // POP RAX
    mem[16'h0C40] = 8'h00;
    mem[16'h0C41] = 8'h81; // ADDN RSP 8
    mem[16'h0C42] = 8'h06;
    mem[16'h0C43] = 8'h08;
    mem[16'h0C44] = 8'h00;
    mem[16'h0C45] = 8'h00;
    mem[16'h0C46] = 8'h00;
    mem[16'h0C47] = 8'h80; // ADD RAX RDI
    mem[16'h0C48] = 8'h00;
    mem[16'h0C49] = 8'h01;
    mem[16'h0C4A] = 8'h85; // SUBN RSP 8
    mem[16'h0C4B] = 8'h06;
    mem[16'h0C4C] = 8'h08;
    mem[16'h0C4D] = 8'h00;
    mem[16'h0C4E] = 8'h00;
    mem[16'h0C4F] = 8'h00;
    mem[16'h0C50] = 8'h04; // PUSH RAX
    mem[16'h0C51] = 8'h00;
    mem[16'h0C52] = 8'h08; // POP RDI
    mem[16'h0C53] = 8'h01;
    mem[16'h0C54] = 8'h81; // ADDN RSP 8
    mem[16'h0C55] = 8'h06;
    mem[16'h0C56] = 8'h08;
    mem[16'h0C57] = 8'h00;
    mem[16'h0C58] = 8'h00;
    mem[16'h0C59] = 8'h00;
    mem[16'h0C5A] = 8'h08; // POP RAX
    mem[16'h0C5B] = 8'h00;
    mem[16'h0C5C] = 8'h81; // ADDN RSP 8
    mem[16'h0C5D] = 8'h06;
    mem[16'h0C5E] = 8'h08;
    mem[16'h0C5F] = 8'h00;
    mem[16'h0C60] = 8'h00;
    mem[16'h0C61] = 8'h00;
    mem[16'h0C62] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0C63] = 8'h00;
    mem[16'h0C64] = 8'h01;
    mem[16'h0C65] = 8'h85; // SUBN RSP 8
    mem[16'h0C66] = 8'h06;
    mem[16'h0C67] = 8'h08;
    mem[16'h0C68] = 8'h00;
    mem[16'h0C69] = 8'h00;
    mem[16'h0C6A] = 8'h00;
    mem[16'h0C6B] = 8'h04; // PUSH RDI
    mem[16'h0C6C] = 8'h01;
    mem[16'h0C6D] = 8'h81; // ADDN RSP 8
    mem[16'h0C6E] = 8'h06;
    mem[16'h0C6F] = 8'h08;
    mem[16'h0C70] = 8'h00;
    mem[16'h0C71] = 8'h00;
    mem[16'h0C72] = 8'h00;
    mem[16'h0C73] = 8'h22; // JMP .Lbegin4
    mem[16'h0C74] = 8'h3F;
    mem[16'h0C75] = 8'h07;
    mem[16'h0C76] = 8'h00;
    mem[16'h0C77] = 8'h00;
    mem[16'h0C78] = 8'h00;
    mem[16'h0C79] = 8'h00;
    mem[16'h0C7A] = 8'h00;
    mem[16'h0C7B] = 8'h00;
                          // .Lend4:
    mem[16'h0C7C] = 8'h85; // SUBN RSP 8
    mem[16'h0C7D] = 8'h06;
    mem[16'h0C7E] = 8'h08;
    mem[16'h0C7F] = 8'h00;
    mem[16'h0C80] = 8'h00;
    mem[16'h0C81] = 8'h00;
    mem[16'h0C82] = 8'h05; // PUSHN 7
    mem[16'h0C83] = 8'h00;
    mem[16'h0C84] = 8'h07;
    mem[16'h0C85] = 8'h00;
    mem[16'h0C86] = 8'h00;
    mem[16'h0C87] = 8'h00;
    mem[16'h0C88] = 8'h40; // MOV RAX RBP
    mem[16'h0C89] = 8'h00;
    mem[16'h0C8A] = 8'h05;
    mem[16'h0C8B] = 8'h85; // SUBN RAX 28
    mem[16'h0C8C] = 8'h00;
    mem[16'h0C8D] = 8'h1C;
    mem[16'h0C8E] = 8'h00;
    mem[16'h0C8F] = 8'h00;
    mem[16'h0C90] = 8'h00;
    mem[16'h0C91] = 8'h85; // SUBN RSP 8
    mem[16'h0C92] = 8'h06;
    mem[16'h0C93] = 8'h08;
    mem[16'h0C94] = 8'h00;
    mem[16'h0C95] = 8'h00;
    mem[16'h0C96] = 8'h00;
    mem[16'h0C97] = 8'h04; // PUSH RAX
    mem[16'h0C98] = 8'h00;
    mem[16'h0C99] = 8'h08; // POP RAX
    mem[16'h0C9A] = 8'h00;
    mem[16'h0C9B] = 8'h81; // ADDN RSP 8
    mem[16'h0C9C] = 8'h06;
    mem[16'h0C9D] = 8'h08;
    mem[16'h0C9E] = 8'h00;
    mem[16'h0C9F] = 8'h00;
    mem[16'h0CA0] = 8'h00;
    mem[16'h0CA1] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0CA2] = 8'h00;
    mem[16'h0CA3] = 8'h00;
    mem[16'h0CA4] = 8'h85; // SUBN RSP 8
    mem[16'h0CA5] = 8'h06;
    mem[16'h0CA6] = 8'h08;
    mem[16'h0CA7] = 8'h00;
    mem[16'h0CA8] = 8'h00;
    mem[16'h0CA9] = 8'h00;
    mem[16'h0CAA] = 8'h04; // PUSH RAX
    mem[16'h0CAB] = 8'h00;
    mem[16'h0CAC] = 8'h08; // POP RDI
    mem[16'h0CAD] = 8'h01;
    mem[16'h0CAE] = 8'h81; // ADDN RSP 8
    mem[16'h0CAF] = 8'h06;
    mem[16'h0CB0] = 8'h08;
    mem[16'h0CB1] = 8'h00;
    mem[16'h0CB2] = 8'h00;
    mem[16'h0CB3] = 8'h00;
    mem[16'h0CB4] = 8'h08; // POP RAX
    mem[16'h0CB5] = 8'h00;
    mem[16'h0CB6] = 8'h81; // ADDN RSP 8
    mem[16'h0CB7] = 8'h06;
    mem[16'h0CB8] = 8'h08;
    mem[16'h0CB9] = 8'h00;
    mem[16'h0CBA] = 8'h00;
    mem[16'h0CBB] = 8'h00;
    mem[16'h0CBC] = 8'h84; // SUB RAX RDI
    mem[16'h0CBD] = 8'h00;
    mem[16'h0CBE] = 8'h01;
    mem[16'h0CBF] = 8'h85; // SUBN RSP 8
    mem[16'h0CC0] = 8'h06;
    mem[16'h0CC1] = 8'h08;
    mem[16'h0CC2] = 8'h00;
    mem[16'h0CC3] = 8'h00;
    mem[16'h0CC4] = 8'h00;
    mem[16'h0CC5] = 8'h04; // PUSH RAX
    mem[16'h0CC6] = 8'h00;
    mem[16'h0CC7] = 8'h40; // MOV RAX RBP
    mem[16'h0CC8] = 8'h00;
    mem[16'h0CC9] = 8'h05;
    mem[16'h0CCA] = 8'h85; // SUBN RAX 32
    mem[16'h0CCB] = 8'h00;
    mem[16'h0CCC] = 8'h20;
    mem[16'h0CCD] = 8'h00;
    mem[16'h0CCE] = 8'h00;
    mem[16'h0CCF] = 8'h00;
    mem[16'h0CD0] = 8'h85; // SUBN RSP 8
    mem[16'h0CD1] = 8'h06;
    mem[16'h0CD2] = 8'h08;
    mem[16'h0CD3] = 8'h00;
    mem[16'h0CD4] = 8'h00;
    mem[16'h0CD5] = 8'h00;
    mem[16'h0CD6] = 8'h04; // PUSH RAX
    mem[16'h0CD7] = 8'h00;
    mem[16'h0CD8] = 8'h08; // POP RAX
    mem[16'h0CD9] = 8'h00;
    mem[16'h0CDA] = 8'h81; // ADDN RSP 8
    mem[16'h0CDB] = 8'h06;
    mem[16'h0CDC] = 8'h08;
    mem[16'h0CDD] = 8'h00;
    mem[16'h0CDE] = 8'h00;
    mem[16'h0CDF] = 8'h00;
    mem[16'h0CE0] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0CE1] = 8'h00;
    mem[16'h0CE2] = 8'h00;
    mem[16'h0CE3] = 8'h85; // SUBN RSP 8
    mem[16'h0CE4] = 8'h06;
    mem[16'h0CE5] = 8'h08;
    mem[16'h0CE6] = 8'h00;
    mem[16'h0CE7] = 8'h00;
    mem[16'h0CE8] = 8'h00;
    mem[16'h0CE9] = 8'h04; // PUSH RAX
    mem[16'h0CEA] = 8'h00;
    mem[16'h0CEB] = 8'h08; // POP RDI
    mem[16'h0CEC] = 8'h01;
    mem[16'h0CED] = 8'h81; // ADDN RSP 8
    mem[16'h0CEE] = 8'h06;
    mem[16'h0CEF] = 8'h08;
    mem[16'h0CF0] = 8'h00;
    mem[16'h0CF1] = 8'h00;
    mem[16'h0CF2] = 8'h00;
    mem[16'h0CF3] = 8'h08; // POP RAX
    mem[16'h0CF4] = 8'h00;
    mem[16'h0CF5] = 8'h81; // ADDN RSP 8
    mem[16'h0CF6] = 8'h06;
    mem[16'h0CF7] = 8'h08;
    mem[16'h0CF8] = 8'h00;
    mem[16'h0CF9] = 8'h00;
    mem[16'h0CFA] = 8'h00;
    mem[16'h0CFB] = 8'h90; // CMP RAX RDI
    mem[16'h0CFC] = 8'h00;
    mem[16'h0CFD] = 8'h01;
    mem[16'h0CFE] = 8'h18; // SETL RAX
    mem[16'h0CFF] = 8'h00;
    mem[16'h0D00] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h0D01] = 8'h00;
    mem[16'h0D02] = 8'h00;
    mem[16'h0D03] = 8'h85; // SUBN RSP 8
    mem[16'h0D04] = 8'h06;
    mem[16'h0D05] = 8'h08;
    mem[16'h0D06] = 8'h00;
    mem[16'h0D07] = 8'h00;
    mem[16'h0D08] = 8'h00;
    mem[16'h0D09] = 8'h04; // PUSH RAX
    mem[16'h0D0A] = 8'h00;
    mem[16'h0D0B] = 8'h08; // POP RAX
    mem[16'h0D0C] = 8'h00;
    mem[16'h0D0D] = 8'h81; // ADDN RSP 8
    mem[16'h0D0E] = 8'h06;
    mem[16'h0D0F] = 8'h08;
    mem[16'h0D10] = 8'h00;
    mem[16'h0D11] = 8'h00;
    mem[16'h0D12] = 8'h00;
    mem[16'h0D13] = 8'h91; // CMPN RAX 0
    mem[16'h0D14] = 8'h00;
    mem[16'h0D15] = 8'h00;
    mem[16'h0D16] = 8'h00;
    mem[16'h0D17] = 8'h00;
    mem[16'h0D18] = 8'h00;
    mem[16'h0D19] = 8'h26; // JE .Lelse8
    mem[16'h0D1A] = 8'hE1;
    mem[16'h0D1B] = 8'h0E;
    mem[16'h0D1C] = 8'h00;
    mem[16'h0D1D] = 8'h00;
    mem[16'h0D1E] = 8'h00;
    mem[16'h0D1F] = 8'h00;
    mem[16'h0D20] = 8'h00;
    mem[16'h0D21] = 8'h00;
    mem[16'h0D22] = 8'h40; // MOV RAX RBP
    mem[16'h0D23] = 8'h00;
    mem[16'h0D24] = 8'h05;
    mem[16'h0D25] = 8'h85; // SUBN RAX 16
    mem[16'h0D26] = 8'h00;
    mem[16'h0D27] = 8'h10;
    mem[16'h0D28] = 8'h00;
    mem[16'h0D29] = 8'h00;
    mem[16'h0D2A] = 8'h00;
    mem[16'h0D2B] = 8'h85; // SUBN RSP 8
    mem[16'h0D2C] = 8'h06;
    mem[16'h0D2D] = 8'h08;
    mem[16'h0D2E] = 8'h00;
    mem[16'h0D2F] = 8'h00;
    mem[16'h0D30] = 8'h00;
    mem[16'h0D31] = 8'h04; // PUSH RAX
    mem[16'h0D32] = 8'h00;
    mem[16'h0D33] = 8'h40; // MOV RAX RBP
    mem[16'h0D34] = 8'h00;
    mem[16'h0D35] = 8'h05;
    mem[16'h0D36] = 8'h85; // SUBN RAX 32
    mem[16'h0D37] = 8'h00;
    mem[16'h0D38] = 8'h20;
    mem[16'h0D39] = 8'h00;
    mem[16'h0D3A] = 8'h00;
    mem[16'h0D3B] = 8'h00;
    mem[16'h0D3C] = 8'h85; // SUBN RSP 8
    mem[16'h0D3D] = 8'h06;
    mem[16'h0D3E] = 8'h08;
    mem[16'h0D3F] = 8'h00;
    mem[16'h0D40] = 8'h00;
    mem[16'h0D41] = 8'h00;
    mem[16'h0D42] = 8'h04; // PUSH RAX
    mem[16'h0D43] = 8'h00;
    mem[16'h0D44] = 8'h08; // POP RAX
    mem[16'h0D45] = 8'h00;
    mem[16'h0D46] = 8'h81; // ADDN RSP 8
    mem[16'h0D47] = 8'h06;
    mem[16'h0D48] = 8'h08;
    mem[16'h0D49] = 8'h00;
    mem[16'h0D4A] = 8'h00;
    mem[16'h0D4B] = 8'h00;
    mem[16'h0D4C] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0D4D] = 8'h00;
    mem[16'h0D4E] = 8'h00;
    mem[16'h0D4F] = 8'h85; // SUBN RSP 8
    mem[16'h0D50] = 8'h06;
    mem[16'h0D51] = 8'h08;
    mem[16'h0D52] = 8'h00;
    mem[16'h0D53] = 8'h00;
    mem[16'h0D54] = 8'h00;
    mem[16'h0D55] = 8'h04; // PUSH RAX
    mem[16'h0D56] = 8'h00;
    mem[16'h0D57] = 8'h40; // MOV RAX RBP
    mem[16'h0D58] = 8'h00;
    mem[16'h0D59] = 8'h05;
    mem[16'h0D5A] = 8'h85; // SUBN RAX 28
    mem[16'h0D5B] = 8'h00;
    mem[16'h0D5C] = 8'h1C;
    mem[16'h0D5D] = 8'h00;
    mem[16'h0D5E] = 8'h00;
    mem[16'h0D5F] = 8'h00;
    mem[16'h0D60] = 8'h85; // SUBN RSP 8
    mem[16'h0D61] = 8'h06;
    mem[16'h0D62] = 8'h08;
    mem[16'h0D63] = 8'h00;
    mem[16'h0D64] = 8'h00;
    mem[16'h0D65] = 8'h00;
    mem[16'h0D66] = 8'h04; // PUSH RAX
    mem[16'h0D67] = 8'h00;
    mem[16'h0D68] = 8'h08; // POP RAX
    mem[16'h0D69] = 8'h00;
    mem[16'h0D6A] = 8'h81; // ADDN RSP 8
    mem[16'h0D6B] = 8'h06;
    mem[16'h0D6C] = 8'h08;
    mem[16'h0D6D] = 8'h00;
    mem[16'h0D6E] = 8'h00;
    mem[16'h0D6F] = 8'h00;
    mem[16'h0D70] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0D71] = 8'h00;
    mem[16'h0D72] = 8'h00;
    mem[16'h0D73] = 8'h85; // SUBN RSP 8
    mem[16'h0D74] = 8'h06;
    mem[16'h0D75] = 8'h08;
    mem[16'h0D76] = 8'h00;
    mem[16'h0D77] = 8'h00;
    mem[16'h0D78] = 8'h00;
    mem[16'h0D79] = 8'h04; // PUSH RAX
    mem[16'h0D7A] = 8'h00;
    mem[16'h0D7B] = 8'h08; // POP RDI
    mem[16'h0D7C] = 8'h01;
    mem[16'h0D7D] = 8'h81; // ADDN RSP 8
    mem[16'h0D7E] = 8'h06;
    mem[16'h0D7F] = 8'h08;
    mem[16'h0D80] = 8'h00;
    mem[16'h0D81] = 8'h00;
    mem[16'h0D82] = 8'h00;
    mem[16'h0D83] = 8'h08; // POP RAX
    mem[16'h0D84] = 8'h00;
    mem[16'h0D85] = 8'h81; // ADDN RSP 8
    mem[16'h0D86] = 8'h06;
    mem[16'h0D87] = 8'h08;
    mem[16'h0D88] = 8'h00;
    mem[16'h0D89] = 8'h00;
    mem[16'h0D8A] = 8'h00;
    mem[16'h0D8B] = 8'h80; // ADD RAX RDI
    mem[16'h0D8C] = 8'h00;
    mem[16'h0D8D] = 8'h01;
    mem[16'h0D8E] = 8'h85; // SUBN RSP 8
    mem[16'h0D8F] = 8'h06;
    mem[16'h0D90] = 8'h08;
    mem[16'h0D91] = 8'h00;
    mem[16'h0D92] = 8'h00;
    mem[16'h0D93] = 8'h00;
    mem[16'h0D94] = 8'h04; // PUSH RAX
    mem[16'h0D95] = 8'h00;
    mem[16'h0D96] = 8'h85; // SUBN RSP 8
    mem[16'h0D97] = 8'h06;
    mem[16'h0D98] = 8'h08;
    mem[16'h0D99] = 8'h00;
    mem[16'h0D9A] = 8'h00;
    mem[16'h0D9B] = 8'h00;
    mem[16'h0D9C] = 8'h05; // PUSHN 7
    mem[16'h0D9D] = 8'h00;
    mem[16'h0D9E] = 8'h07;
    mem[16'h0D9F] = 8'h00;
    mem[16'h0DA0] = 8'h00;
    mem[16'h0DA1] = 8'h00;
    mem[16'h0DA2] = 8'h08; // POP RDI
    mem[16'h0DA3] = 8'h01;
    mem[16'h0DA4] = 8'h81; // ADDN RSP 8
    mem[16'h0DA5] = 8'h06;
    mem[16'h0DA6] = 8'h08;
    mem[16'h0DA7] = 8'h00;
    mem[16'h0DA8] = 8'h00;
    mem[16'h0DA9] = 8'h00;
    mem[16'h0DAA] = 8'h08; // POP RAX
    mem[16'h0DAB] = 8'h00;
    mem[16'h0DAC] = 8'h81; // ADDN RSP 8
    mem[16'h0DAD] = 8'h06;
    mem[16'h0DAE] = 8'h08;
    mem[16'h0DAF] = 8'h00;
    mem[16'h0DB0] = 8'h00;
    mem[16'h0DB1] = 8'h00;
    mem[16'h0DB2] = 8'h84; // SUB RAX RDI
    mem[16'h0DB3] = 8'h00;
    mem[16'h0DB4] = 8'h01;
    mem[16'h0DB5] = 8'h85; // SUBN RSP 8
    mem[16'h0DB6] = 8'h06;
    mem[16'h0DB7] = 8'h08;
    mem[16'h0DB8] = 8'h00;
    mem[16'h0DB9] = 8'h00;
    mem[16'h0DBA] = 8'h00;
    mem[16'h0DBB] = 8'h04; // PUSH RAX
    mem[16'h0DBC] = 8'h00;
    mem[16'h0DBD] = 8'h08; // POP RDI
    mem[16'h0DBE] = 8'h01;
    mem[16'h0DBF] = 8'h81; // ADDN RSP 8
    mem[16'h0DC0] = 8'h06;
    mem[16'h0DC1] = 8'h08;
    mem[16'h0DC2] = 8'h00;
    mem[16'h0DC3] = 8'h00;
    mem[16'h0DC4] = 8'h00;
    mem[16'h0DC5] = 8'h08; // POP RAX
    mem[16'h0DC6] = 8'h00;
    mem[16'h0DC7] = 8'h81; // ADDN RSP 8
    mem[16'h0DC8] = 8'h06;
    mem[16'h0DC9] = 8'h08;
    mem[16'h0DCA] = 8'h00;
    mem[16'h0DCB] = 8'h00;
    mem[16'h0DCC] = 8'h00;
    mem[16'h0DCD] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0DCE] = 8'h00;
    mem[16'h0DCF] = 8'h01;
    mem[16'h0DD0] = 8'h85; // SUBN RSP 8
    mem[16'h0DD1] = 8'h06;
    mem[16'h0DD2] = 8'h08;
    mem[16'h0DD3] = 8'h00;
    mem[16'h0DD4] = 8'h00;
    mem[16'h0DD5] = 8'h00;
    mem[16'h0DD6] = 8'h04; // PUSH RDI
    mem[16'h0DD7] = 8'h01;
    mem[16'h0DD8] = 8'h81; // ADDN RSP 8
    mem[16'h0DD9] = 8'h06;
    mem[16'h0DDA] = 8'h08;
    mem[16'h0DDB] = 8'h00;
    mem[16'h0DDC] = 8'h00;
    mem[16'h0DDD] = 8'h00;
    mem[16'h0DDE] = 8'h40; // MOV RAX RBP
    mem[16'h0DDF] = 8'h00;
    mem[16'h0DE0] = 8'h05;
    mem[16'h0DE1] = 8'h85; // SUBN RAX 12
    mem[16'h0DE2] = 8'h00;
    mem[16'h0DE3] = 8'h0C;
    mem[16'h0DE4] = 8'h00;
    mem[16'h0DE5] = 8'h00;
    mem[16'h0DE6] = 8'h00;
    mem[16'h0DE7] = 8'h85; // SUBN RSP 8
    mem[16'h0DE8] = 8'h06;
    mem[16'h0DE9] = 8'h08;
    mem[16'h0DEA] = 8'h00;
    mem[16'h0DEB] = 8'h00;
    mem[16'h0DEC] = 8'h00;
    mem[16'h0DED] = 8'h04; // PUSH RAX
    mem[16'h0DEE] = 8'h00;
    mem[16'h0DEF] = 8'h85; // SUBN RSP 8
    mem[16'h0DF0] = 8'h06;
    mem[16'h0DF1] = 8'h08;
    mem[16'h0DF2] = 8'h00;
    mem[16'h0DF3] = 8'h00;
    mem[16'h0DF4] = 8'h00;
    mem[16'h0DF5] = 8'h05; // PUSHN 7
    mem[16'h0DF6] = 8'h00;
    mem[16'h0DF7] = 8'h07;
    mem[16'h0DF8] = 8'h00;
    mem[16'h0DF9] = 8'h00;
    mem[16'h0DFA] = 8'h00;
    mem[16'h0DFB] = 8'h08; // POP RDI
    mem[16'h0DFC] = 8'h01;
    mem[16'h0DFD] = 8'h81; // ADDN RSP 8
    mem[16'h0DFE] = 8'h06;
    mem[16'h0DFF] = 8'h08;
    mem[16'h0E00] = 8'h00;
    mem[16'h0E01] = 8'h00;
    mem[16'h0E02] = 8'h00;
    mem[16'h0E03] = 8'h08; // POP RAX
    mem[16'h0E04] = 8'h00;
    mem[16'h0E05] = 8'h81; // ADDN RSP 8
    mem[16'h0E06] = 8'h06;
    mem[16'h0E07] = 8'h08;
    mem[16'h0E08] = 8'h00;
    mem[16'h0E09] = 8'h00;
    mem[16'h0E0A] = 8'h00;
    mem[16'h0E0B] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0E0C] = 8'h00;
    mem[16'h0E0D] = 8'h01;
    mem[16'h0E0E] = 8'h85; // SUBN RSP 8
    mem[16'h0E0F] = 8'h06;
    mem[16'h0E10] = 8'h08;
    mem[16'h0E11] = 8'h00;
    mem[16'h0E12] = 8'h00;
    mem[16'h0E13] = 8'h00;
    mem[16'h0E14] = 8'h04; // PUSH RDI
    mem[16'h0E15] = 8'h01;
    mem[16'h0E16] = 8'h81; // ADDN RSP 8
    mem[16'h0E17] = 8'h06;
    mem[16'h0E18] = 8'h08;
    mem[16'h0E19] = 8'h00;
    mem[16'h0E1A] = 8'h00;
    mem[16'h0E1B] = 8'h00;
    mem[16'h0E1C] = 8'h40; // MOV RAX RBP
    mem[16'h0E1D] = 8'h00;
    mem[16'h0E1E] = 8'h05;
    mem[16'h0E1F] = 8'h85; // SUBN RAX 8
    mem[16'h0E20] = 8'h00;
    mem[16'h0E21] = 8'h08;
    mem[16'h0E22] = 8'h00;
    mem[16'h0E23] = 8'h00;
    mem[16'h0E24] = 8'h00;
    mem[16'h0E25] = 8'h85; // SUBN RSP 8
    mem[16'h0E26] = 8'h06;
    mem[16'h0E27] = 8'h08;
    mem[16'h0E28] = 8'h00;
    mem[16'h0E29] = 8'h00;
    mem[16'h0E2A] = 8'h00;
    mem[16'h0E2B] = 8'h04; // PUSH RAX
    mem[16'h0E2C] = 8'h00;
    mem[16'h0E2D] = 8'h85; // SUBN RSP 8
    mem[16'h0E2E] = 8'h06;
    mem[16'h0E2F] = 8'h08;
    mem[16'h0E30] = 8'h00;
    mem[16'h0E31] = 8'h00;
    mem[16'h0E32] = 8'h00;
    mem[16'h0E33] = 8'h05; // PUSHN 15
    mem[16'h0E34] = 8'h00;
    mem[16'h0E35] = 8'h0F;
    mem[16'h0E36] = 8'h00;
    mem[16'h0E37] = 8'h00;
    mem[16'h0E38] = 8'h00;
    mem[16'h0E39] = 8'h40; // MOV RAX RBP
    mem[16'h0E3A] = 8'h00;
    mem[16'h0E3B] = 8'h05;
    mem[16'h0E3C] = 8'h85; // SUBN RAX 32
    mem[16'h0E3D] = 8'h00;
    mem[16'h0E3E] = 8'h20;
    mem[16'h0E3F] = 8'h00;
    mem[16'h0E40] = 8'h00;
    mem[16'h0E41] = 8'h00;
    mem[16'h0E42] = 8'h85; // SUBN RSP 8
    mem[16'h0E43] = 8'h06;
    mem[16'h0E44] = 8'h08;
    mem[16'h0E45] = 8'h00;
    mem[16'h0E46] = 8'h00;
    mem[16'h0E47] = 8'h00;
    mem[16'h0E48] = 8'h04; // PUSH RAX
    mem[16'h0E49] = 8'h00;
    mem[16'h0E4A] = 8'h08; // POP RAX
    mem[16'h0E4B] = 8'h00;
    mem[16'h0E4C] = 8'h81; // ADDN RSP 8
    mem[16'h0E4D] = 8'h06;
    mem[16'h0E4E] = 8'h08;
    mem[16'h0E4F] = 8'h00;
    mem[16'h0E50] = 8'h00;
    mem[16'h0E51] = 8'h00;
    mem[16'h0E52] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0E53] = 8'h00;
    mem[16'h0E54] = 8'h00;
    mem[16'h0E55] = 8'h85; // SUBN RSP 8
    mem[16'h0E56] = 8'h06;
    mem[16'h0E57] = 8'h08;
    mem[16'h0E58] = 8'h00;
    mem[16'h0E59] = 8'h00;
    mem[16'h0E5A] = 8'h00;
    mem[16'h0E5B] = 8'h04; // PUSH RAX
    mem[16'h0E5C] = 8'h00;
    mem[16'h0E5D] = 8'h40; // MOV RAX RBP
    mem[16'h0E5E] = 8'h00;
    mem[16'h0E5F] = 8'h05;
    mem[16'h0E60] = 8'h85; // SUBN RAX 28
    mem[16'h0E61] = 8'h00;
    mem[16'h0E62] = 8'h1C;
    mem[16'h0E63] = 8'h00;
    mem[16'h0E64] = 8'h00;
    mem[16'h0E65] = 8'h00;
    mem[16'h0E66] = 8'h85; // SUBN RSP 8
    mem[16'h0E67] = 8'h06;
    mem[16'h0E68] = 8'h08;
    mem[16'h0E69] = 8'h00;
    mem[16'h0E6A] = 8'h00;
    mem[16'h0E6B] = 8'h00;
    mem[16'h0E6C] = 8'h04; // PUSH RAX
    mem[16'h0E6D] = 8'h00;
    mem[16'h0E6E] = 8'h08; // POP RAX
    mem[16'h0E6F] = 8'h00;
    mem[16'h0E70] = 8'h81; // ADDN RSP 8
    mem[16'h0E71] = 8'h06;
    mem[16'h0E72] = 8'h08;
    mem[16'h0E73] = 8'h00;
    mem[16'h0E74] = 8'h00;
    mem[16'h0E75] = 8'h00;
    mem[16'h0E76] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0E77] = 8'h00;
    mem[16'h0E78] = 8'h00;
    mem[16'h0E79] = 8'h85; // SUBN RSP 8
    mem[16'h0E7A] = 8'h06;
    mem[16'h0E7B] = 8'h08;
    mem[16'h0E7C] = 8'h00;
    mem[16'h0E7D] = 8'h00;
    mem[16'h0E7E] = 8'h00;
    mem[16'h0E7F] = 8'h04; // PUSH RAX
    mem[16'h0E80] = 8'h00;
    mem[16'h0E81] = 8'h08; // POP RDI
    mem[16'h0E82] = 8'h01;
    mem[16'h0E83] = 8'h81; // ADDN RSP 8
    mem[16'h0E84] = 8'h06;
    mem[16'h0E85] = 8'h08;
    mem[16'h0E86] = 8'h00;
    mem[16'h0E87] = 8'h00;
    mem[16'h0E88] = 8'h00;
    mem[16'h0E89] = 8'h08; // POP RAX
    mem[16'h0E8A] = 8'h00;
    mem[16'h0E8B] = 8'h81; // ADDN RSP 8
    mem[16'h0E8C] = 8'h06;
    mem[16'h0E8D] = 8'h08;
    mem[16'h0E8E] = 8'h00;
    mem[16'h0E8F] = 8'h00;
    mem[16'h0E90] = 8'h00;
    mem[16'h0E91] = 8'h80; // ADD RAX RDI
    mem[16'h0E92] = 8'h00;
    mem[16'h0E93] = 8'h01;
    mem[16'h0E94] = 8'h85; // SUBN RSP 8
    mem[16'h0E95] = 8'h06;
    mem[16'h0E96] = 8'h08;
    mem[16'h0E97] = 8'h00;
    mem[16'h0E98] = 8'h00;
    mem[16'h0E99] = 8'h00;
    mem[16'h0E9A] = 8'h04; // PUSH RAX
    mem[16'h0E9B] = 8'h00;
    mem[16'h0E9C] = 8'h08; // POP RDI
    mem[16'h0E9D] = 8'h01;
    mem[16'h0E9E] = 8'h81; // ADDN RSP 8
    mem[16'h0E9F] = 8'h06;
    mem[16'h0EA0] = 8'h08;
    mem[16'h0EA1] = 8'h00;
    mem[16'h0EA2] = 8'h00;
    mem[16'h0EA3] = 8'h00;
    mem[16'h0EA4] = 8'h08; // POP RAX
    mem[16'h0EA5] = 8'h00;
    mem[16'h0EA6] = 8'h81; // ADDN RSP 8
    mem[16'h0EA7] = 8'h06;
    mem[16'h0EA8] = 8'h08;
    mem[16'h0EA9] = 8'h00;
    mem[16'h0EAA] = 8'h00;
    mem[16'h0EAB] = 8'h00;
    mem[16'h0EAC] = 8'h84; // SUB RAX RDI
    mem[16'h0EAD] = 8'h00;
    mem[16'h0EAE] = 8'h01;
    mem[16'h0EAF] = 8'h85; // SUBN RSP 8
    mem[16'h0EB0] = 8'h06;
    mem[16'h0EB1] = 8'h08;
    mem[16'h0EB2] = 8'h00;
    mem[16'h0EB3] = 8'h00;
    mem[16'h0EB4] = 8'h00;
    mem[16'h0EB5] = 8'h04; // PUSH RAX
    mem[16'h0EB6] = 8'h00;
    mem[16'h0EB7] = 8'h08; // POP RDI
    mem[16'h0EB8] = 8'h01;
    mem[16'h0EB9] = 8'h81; // ADDN RSP 8
    mem[16'h0EBA] = 8'h06;
    mem[16'h0EBB] = 8'h08;
    mem[16'h0EBC] = 8'h00;
    mem[16'h0EBD] = 8'h00;
    mem[16'h0EBE] = 8'h00;
    mem[16'h0EBF] = 8'h08; // POP RAX
    mem[16'h0EC0] = 8'h00;
    mem[16'h0EC1] = 8'h81; // ADDN RSP 8
    mem[16'h0EC2] = 8'h06;
    mem[16'h0EC3] = 8'h08;
    mem[16'h0EC4] = 8'h00;
    mem[16'h0EC5] = 8'h00;
    mem[16'h0EC6] = 8'h00;
    mem[16'h0EC7] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0EC8] = 8'h00;
    mem[16'h0EC9] = 8'h01;
    mem[16'h0ECA] = 8'h85; // SUBN RSP 8
    mem[16'h0ECB] = 8'h06;
    mem[16'h0ECC] = 8'h08;
    mem[16'h0ECD] = 8'h00;
    mem[16'h0ECE] = 8'h00;
    mem[16'h0ECF] = 8'h00;
    mem[16'h0ED0] = 8'h04; // PUSH RDI
    mem[16'h0ED1] = 8'h01;
    mem[16'h0ED2] = 8'h81; // ADDN RSP 8
    mem[16'h0ED3] = 8'h06;
    mem[16'h0ED4] = 8'h08;
    mem[16'h0ED5] = 8'h00;
    mem[16'h0ED6] = 8'h00;
    mem[16'h0ED7] = 8'h00;
    mem[16'h0ED8] = 8'h22; // JMP .Lend8
    mem[16'h0ED9] = 8'h70;
    mem[16'h0EDA] = 8'h10;
    mem[16'h0EDB] = 8'h00;
    mem[16'h0EDC] = 8'h00;
    mem[16'h0EDD] = 8'h00;
    mem[16'h0EDE] = 8'h00;
    mem[16'h0EDF] = 8'h00;
    mem[16'h0EE0] = 8'h00;
                          // .Lelse8:
    mem[16'h0EE1] = 8'h40; // MOV RAX RBP
    mem[16'h0EE2] = 8'h00;
    mem[16'h0EE3] = 8'h05;
    mem[16'h0EE4] = 8'h85; // SUBN RAX 16
    mem[16'h0EE5] = 8'h00;
    mem[16'h0EE6] = 8'h10;
    mem[16'h0EE7] = 8'h00;
    mem[16'h0EE8] = 8'h00;
    mem[16'h0EE9] = 8'h00;
    mem[16'h0EEA] = 8'h85; // SUBN RSP 8
    mem[16'h0EEB] = 8'h06;
    mem[16'h0EEC] = 8'h08;
    mem[16'h0EED] = 8'h00;
    mem[16'h0EEE] = 8'h00;
    mem[16'h0EEF] = 8'h00;
    mem[16'h0EF0] = 8'h04; // PUSH RAX
    mem[16'h0EF1] = 8'h00;
    mem[16'h0EF2] = 8'h85; // SUBN RSP 8
    mem[16'h0EF3] = 8'h06;
    mem[16'h0EF4] = 8'h08;
    mem[16'h0EF5] = 8'h00;
    mem[16'h0EF6] = 8'h00;
    mem[16'h0EF7] = 8'h00;
    mem[16'h0EF8] = 8'h05; // PUSHN 0
    mem[16'h0EF9] = 8'h00;
    mem[16'h0EFA] = 8'h00;
    mem[16'h0EFB] = 8'h00;
    mem[16'h0EFC] = 8'h00;
    mem[16'h0EFD] = 8'h00;
    mem[16'h0EFE] = 8'h08; // POP RDI
    mem[16'h0EFF] = 8'h01;
    mem[16'h0F00] = 8'h81; // ADDN RSP 8
    mem[16'h0F01] = 8'h06;
    mem[16'h0F02] = 8'h08;
    mem[16'h0F03] = 8'h00;
    mem[16'h0F04] = 8'h00;
    mem[16'h0F05] = 8'h00;
    mem[16'h0F06] = 8'h08; // POP RAX
    mem[16'h0F07] = 8'h00;
    mem[16'h0F08] = 8'h81; // ADDN RSP 8
    mem[16'h0F09] = 8'h06;
    mem[16'h0F0A] = 8'h08;
    mem[16'h0F0B] = 8'h00;
    mem[16'h0F0C] = 8'h00;
    mem[16'h0F0D] = 8'h00;
    mem[16'h0F0E] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0F0F] = 8'h00;
    mem[16'h0F10] = 8'h01;
    mem[16'h0F11] = 8'h85; // SUBN RSP 8
    mem[16'h0F12] = 8'h06;
    mem[16'h0F13] = 8'h08;
    mem[16'h0F14] = 8'h00;
    mem[16'h0F15] = 8'h00;
    mem[16'h0F16] = 8'h00;
    mem[16'h0F17] = 8'h04; // PUSH RDI
    mem[16'h0F18] = 8'h01;
    mem[16'h0F19] = 8'h81; // ADDN RSP 8
    mem[16'h0F1A] = 8'h06;
    mem[16'h0F1B] = 8'h08;
    mem[16'h0F1C] = 8'h00;
    mem[16'h0F1D] = 8'h00;
    mem[16'h0F1E] = 8'h00;
    mem[16'h0F1F] = 8'h40; // MOV RAX RBP
    mem[16'h0F20] = 8'h00;
    mem[16'h0F21] = 8'h05;
    mem[16'h0F22] = 8'h85; // SUBN RAX 12
    mem[16'h0F23] = 8'h00;
    mem[16'h0F24] = 8'h0C;
    mem[16'h0F25] = 8'h00;
    mem[16'h0F26] = 8'h00;
    mem[16'h0F27] = 8'h00;
    mem[16'h0F28] = 8'h85; // SUBN RSP 8
    mem[16'h0F29] = 8'h06;
    mem[16'h0F2A] = 8'h08;
    mem[16'h0F2B] = 8'h00;
    mem[16'h0F2C] = 8'h00;
    mem[16'h0F2D] = 8'h00;
    mem[16'h0F2E] = 8'h04; // PUSH RAX
    mem[16'h0F2F] = 8'h00;
    mem[16'h0F30] = 8'h40; // MOV RAX RBP
    mem[16'h0F31] = 8'h00;
    mem[16'h0F32] = 8'h05;
    mem[16'h0F33] = 8'h85; // SUBN RAX 32
    mem[16'h0F34] = 8'h00;
    mem[16'h0F35] = 8'h20;
    mem[16'h0F36] = 8'h00;
    mem[16'h0F37] = 8'h00;
    mem[16'h0F38] = 8'h00;
    mem[16'h0F39] = 8'h85; // SUBN RSP 8
    mem[16'h0F3A] = 8'h06;
    mem[16'h0F3B] = 8'h08;
    mem[16'h0F3C] = 8'h00;
    mem[16'h0F3D] = 8'h00;
    mem[16'h0F3E] = 8'h00;
    mem[16'h0F3F] = 8'h04; // PUSH RAX
    mem[16'h0F40] = 8'h00;
    mem[16'h0F41] = 8'h08; // POP RAX
    mem[16'h0F42] = 8'h00;
    mem[16'h0F43] = 8'h81; // ADDN RSP 8
    mem[16'h0F44] = 8'h06;
    mem[16'h0F45] = 8'h08;
    mem[16'h0F46] = 8'h00;
    mem[16'h0F47] = 8'h00;
    mem[16'h0F48] = 8'h00;
    mem[16'h0F49] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0F4A] = 8'h00;
    mem[16'h0F4B] = 8'h00;
    mem[16'h0F4C] = 8'h85; // SUBN RSP 8
    mem[16'h0F4D] = 8'h06;
    mem[16'h0F4E] = 8'h08;
    mem[16'h0F4F] = 8'h00;
    mem[16'h0F50] = 8'h00;
    mem[16'h0F51] = 8'h00;
    mem[16'h0F52] = 8'h04; // PUSH RAX
    mem[16'h0F53] = 8'h00;
    mem[16'h0F54] = 8'h40; // MOV RAX RBP
    mem[16'h0F55] = 8'h00;
    mem[16'h0F56] = 8'h05;
    mem[16'h0F57] = 8'h85; // SUBN RAX 28
    mem[16'h0F58] = 8'h00;
    mem[16'h0F59] = 8'h1C;
    mem[16'h0F5A] = 8'h00;
    mem[16'h0F5B] = 8'h00;
    mem[16'h0F5C] = 8'h00;
    mem[16'h0F5D] = 8'h85; // SUBN RSP 8
    mem[16'h0F5E] = 8'h06;
    mem[16'h0F5F] = 8'h08;
    mem[16'h0F60] = 8'h00;
    mem[16'h0F61] = 8'h00;
    mem[16'h0F62] = 8'h00;
    mem[16'h0F63] = 8'h04; // PUSH RAX
    mem[16'h0F64] = 8'h00;
    mem[16'h0F65] = 8'h08; // POP RAX
    mem[16'h0F66] = 8'h00;
    mem[16'h0F67] = 8'h81; // ADDN RSP 8
    mem[16'h0F68] = 8'h06;
    mem[16'h0F69] = 8'h08;
    mem[16'h0F6A] = 8'h00;
    mem[16'h0F6B] = 8'h00;
    mem[16'h0F6C] = 8'h00;
    mem[16'h0F6D] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0F6E] = 8'h00;
    mem[16'h0F6F] = 8'h00;
    mem[16'h0F70] = 8'h85; // SUBN RSP 8
    mem[16'h0F71] = 8'h06;
    mem[16'h0F72] = 8'h08;
    mem[16'h0F73] = 8'h00;
    mem[16'h0F74] = 8'h00;
    mem[16'h0F75] = 8'h00;
    mem[16'h0F76] = 8'h04; // PUSH RAX
    mem[16'h0F77] = 8'h00;
    mem[16'h0F78] = 8'h08; // POP RDI
    mem[16'h0F79] = 8'h01;
    mem[16'h0F7A] = 8'h81; // ADDN RSP 8
    mem[16'h0F7B] = 8'h06;
    mem[16'h0F7C] = 8'h08;
    mem[16'h0F7D] = 8'h00;
    mem[16'h0F7E] = 8'h00;
    mem[16'h0F7F] = 8'h00;
    mem[16'h0F80] = 8'h08; // POP RAX
    mem[16'h0F81] = 8'h00;
    mem[16'h0F82] = 8'h81; // ADDN RSP 8
    mem[16'h0F83] = 8'h06;
    mem[16'h0F84] = 8'h08;
    mem[16'h0F85] = 8'h00;
    mem[16'h0F86] = 8'h00;
    mem[16'h0F87] = 8'h00;
    mem[16'h0F88] = 8'h80; // ADD RAX RDI
    mem[16'h0F89] = 8'h00;
    mem[16'h0F8A] = 8'h01;
    mem[16'h0F8B] = 8'h85; // SUBN RSP 8
    mem[16'h0F8C] = 8'h06;
    mem[16'h0F8D] = 8'h08;
    mem[16'h0F8E] = 8'h00;
    mem[16'h0F8F] = 8'h00;
    mem[16'h0F90] = 8'h00;
    mem[16'h0F91] = 8'h04; // PUSH RAX
    mem[16'h0F92] = 8'h00;
    mem[16'h0F93] = 8'h08; // POP RDI
    mem[16'h0F94] = 8'h01;
    mem[16'h0F95] = 8'h81; // ADDN RSP 8
    mem[16'h0F96] = 8'h06;
    mem[16'h0F97] = 8'h08;
    mem[16'h0F98] = 8'h00;
    mem[16'h0F99] = 8'h00;
    mem[16'h0F9A] = 8'h00;
    mem[16'h0F9B] = 8'h08; // POP RAX
    mem[16'h0F9C] = 8'h00;
    mem[16'h0F9D] = 8'h81; // ADDN RSP 8
    mem[16'h0F9E] = 8'h06;
    mem[16'h0F9F] = 8'h08;
    mem[16'h0FA0] = 8'h00;
    mem[16'h0FA1] = 8'h00;
    mem[16'h0FA2] = 8'h00;
    mem[16'h0FA3] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h0FA4] = 8'h00;
    mem[16'h0FA5] = 8'h01;
    mem[16'h0FA6] = 8'h85; // SUBN RSP 8
    mem[16'h0FA7] = 8'h06;
    mem[16'h0FA8] = 8'h08;
    mem[16'h0FA9] = 8'h00;
    mem[16'h0FAA] = 8'h00;
    mem[16'h0FAB] = 8'h00;
    mem[16'h0FAC] = 8'h04; // PUSH RDI
    mem[16'h0FAD] = 8'h01;
    mem[16'h0FAE] = 8'h81; // ADDN RSP 8
    mem[16'h0FAF] = 8'h06;
    mem[16'h0FB0] = 8'h08;
    mem[16'h0FB1] = 8'h00;
    mem[16'h0FB2] = 8'h00;
    mem[16'h0FB3] = 8'h00;
    mem[16'h0FB4] = 8'h40; // MOV RAX RBP
    mem[16'h0FB5] = 8'h00;
    mem[16'h0FB6] = 8'h05;
    mem[16'h0FB7] = 8'h85; // SUBN RAX 8
    mem[16'h0FB8] = 8'h00;
    mem[16'h0FB9] = 8'h08;
    mem[16'h0FBA] = 8'h00;
    mem[16'h0FBB] = 8'h00;
    mem[16'h0FBC] = 8'h00;
    mem[16'h0FBD] = 8'h85; // SUBN RSP 8
    mem[16'h0FBE] = 8'h06;
    mem[16'h0FBF] = 8'h08;
    mem[16'h0FC0] = 8'h00;
    mem[16'h0FC1] = 8'h00;
    mem[16'h0FC2] = 8'h00;
    mem[16'h0FC3] = 8'h04; // PUSH RAX
    mem[16'h0FC4] = 8'h00;
    mem[16'h0FC5] = 8'h40; // MOV RAX RBP
    mem[16'h0FC6] = 8'h00;
    mem[16'h0FC7] = 8'h05;
    mem[16'h0FC8] = 8'h85; // SUBN RAX 32
    mem[16'h0FC9] = 8'h00;
    mem[16'h0FCA] = 8'h20;
    mem[16'h0FCB] = 8'h00;
    mem[16'h0FCC] = 8'h00;
    mem[16'h0FCD] = 8'h00;
    mem[16'h0FCE] = 8'h85; // SUBN RSP 8
    mem[16'h0FCF] = 8'h06;
    mem[16'h0FD0] = 8'h08;
    mem[16'h0FD1] = 8'h00;
    mem[16'h0FD2] = 8'h00;
    mem[16'h0FD3] = 8'h00;
    mem[16'h0FD4] = 8'h04; // PUSH RAX
    mem[16'h0FD5] = 8'h00;
    mem[16'h0FD6] = 8'h08; // POP RAX
    mem[16'h0FD7] = 8'h00;
    mem[16'h0FD8] = 8'h81; // ADDN RSP 8
    mem[16'h0FD9] = 8'h06;
    mem[16'h0FDA] = 8'h08;
    mem[16'h0FDB] = 8'h00;
    mem[16'h0FDC] = 8'h00;
    mem[16'h0FDD] = 8'h00;
    mem[16'h0FDE] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h0FDF] = 8'h00;
    mem[16'h0FE0] = 8'h00;
    mem[16'h0FE1] = 8'h85; // SUBN RSP 8
    mem[16'h0FE2] = 8'h06;
    mem[16'h0FE3] = 8'h08;
    mem[16'h0FE4] = 8'h00;
    mem[16'h0FE5] = 8'h00;
    mem[16'h0FE6] = 8'h00;
    mem[16'h0FE7] = 8'h04; // PUSH RAX
    mem[16'h0FE8] = 8'h00;
    mem[16'h0FE9] = 8'h40; // MOV RAX RBP
    mem[16'h0FEA] = 8'h00;
    mem[16'h0FEB] = 8'h05;
    mem[16'h0FEC] = 8'h85; // SUBN RAX 28
    mem[16'h0FED] = 8'h00;
    mem[16'h0FEE] = 8'h1C;
    mem[16'h0FEF] = 8'h00;
    mem[16'h0FF0] = 8'h00;
    mem[16'h0FF1] = 8'h00;
    mem[16'h0FF2] = 8'h85; // SUBN RSP 8
    mem[16'h0FF3] = 8'h06;
    mem[16'h0FF4] = 8'h08;
    mem[16'h0FF5] = 8'h00;
    mem[16'h0FF6] = 8'h00;
    mem[16'h0FF7] = 8'h00;
    mem[16'h0FF8] = 8'h04; // PUSH RAX
    mem[16'h0FF9] = 8'h00;
    mem[16'h0FFA] = 8'h08; // POP RAX
    mem[16'h0FFB] = 8'h00;
    mem[16'h0FFC] = 8'h81; // ADDN RSP 8
    mem[16'h0FFD] = 8'h06;
    mem[16'h0FFE] = 8'h08;
    mem[16'h0FFF] = 8'h00;
    mem[16'h1000] = 8'h00;
    mem[16'h1001] = 8'h00;
    mem[16'h1002] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1003] = 8'h00;
    mem[16'h1004] = 8'h00;
    mem[16'h1005] = 8'h85; // SUBN RSP 8
    mem[16'h1006] = 8'h06;
    mem[16'h1007] = 8'h08;
    mem[16'h1008] = 8'h00;
    mem[16'h1009] = 8'h00;
    mem[16'h100A] = 8'h00;
    mem[16'h100B] = 8'h04; // PUSH RAX
    mem[16'h100C] = 8'h00;
    mem[16'h100D] = 8'h08; // POP RDI
    mem[16'h100E] = 8'h01;
    mem[16'h100F] = 8'h81; // ADDN RSP 8
    mem[16'h1010] = 8'h06;
    mem[16'h1011] = 8'h08;
    mem[16'h1012] = 8'h00;
    mem[16'h1013] = 8'h00;
    mem[16'h1014] = 8'h00;
    mem[16'h1015] = 8'h08; // POP RAX
    mem[16'h1016] = 8'h00;
    mem[16'h1017] = 8'h81; // ADDN RSP 8
    mem[16'h1018] = 8'h06;
    mem[16'h1019] = 8'h08;
    mem[16'h101A] = 8'h00;
    mem[16'h101B] = 8'h00;
    mem[16'h101C] = 8'h00;
    mem[16'h101D] = 8'h80; // ADD RAX RDI
    mem[16'h101E] = 8'h00;
    mem[16'h101F] = 8'h01;
    mem[16'h1020] = 8'h85; // SUBN RSP 8
    mem[16'h1021] = 8'h06;
    mem[16'h1022] = 8'h08;
    mem[16'h1023] = 8'h00;
    mem[16'h1024] = 8'h00;
    mem[16'h1025] = 8'h00;
    mem[16'h1026] = 8'h04; // PUSH RAX
    mem[16'h1027] = 8'h00;
    mem[16'h1028] = 8'h85; // SUBN RSP 8
    mem[16'h1029] = 8'h06;
    mem[16'h102A] = 8'h08;
    mem[16'h102B] = 8'h00;
    mem[16'h102C] = 8'h00;
    mem[16'h102D] = 8'h00;
    mem[16'h102E] = 8'h05; // PUSHN 1
    mem[16'h102F] = 8'h00;
    mem[16'h1030] = 8'h01;
    mem[16'h1031] = 8'h00;
    mem[16'h1032] = 8'h00;
    mem[16'h1033] = 8'h00;
    mem[16'h1034] = 8'h08; // POP RDI
    mem[16'h1035] = 8'h01;
    mem[16'h1036] = 8'h81; // ADDN RSP 8
    mem[16'h1037] = 8'h06;
    mem[16'h1038] = 8'h08;
    mem[16'h1039] = 8'h00;
    mem[16'h103A] = 8'h00;
    mem[16'h103B] = 8'h00;
    mem[16'h103C] = 8'h08; // POP RAX
    mem[16'h103D] = 8'h00;
    mem[16'h103E] = 8'h81; // ADDN RSP 8
    mem[16'h103F] = 8'h06;
    mem[16'h1040] = 8'h08;
    mem[16'h1041] = 8'h00;
    mem[16'h1042] = 8'h00;
    mem[16'h1043] = 8'h00;
    mem[16'h1044] = 8'h80; // ADD RAX RDI
    mem[16'h1045] = 8'h00;
    mem[16'h1046] = 8'h01;
    mem[16'h1047] = 8'h85; // SUBN RSP 8
    mem[16'h1048] = 8'h06;
    mem[16'h1049] = 8'h08;
    mem[16'h104A] = 8'h00;
    mem[16'h104B] = 8'h00;
    mem[16'h104C] = 8'h00;
    mem[16'h104D] = 8'h04; // PUSH RAX
    mem[16'h104E] = 8'h00;
    mem[16'h104F] = 8'h08; // POP RDI
    mem[16'h1050] = 8'h01;
    mem[16'h1051] = 8'h81; // ADDN RSP 8
    mem[16'h1052] = 8'h06;
    mem[16'h1053] = 8'h08;
    mem[16'h1054] = 8'h00;
    mem[16'h1055] = 8'h00;
    mem[16'h1056] = 8'h00;
    mem[16'h1057] = 8'h08; // POP RAX
    mem[16'h1058] = 8'h00;
    mem[16'h1059] = 8'h81; // ADDN RSP 8
    mem[16'h105A] = 8'h06;
    mem[16'h105B] = 8'h08;
    mem[16'h105C] = 8'h00;
    mem[16'h105D] = 8'h00;
    mem[16'h105E] = 8'h00;
    mem[16'h105F] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h1060] = 8'h00;
    mem[16'h1061] = 8'h01;
    mem[16'h1062] = 8'h85; // SUBN RSP 8
    mem[16'h1063] = 8'h06;
    mem[16'h1064] = 8'h08;
    mem[16'h1065] = 8'h00;
    mem[16'h1066] = 8'h00;
    mem[16'h1067] = 8'h00;
    mem[16'h1068] = 8'h04; // PUSH RDI
    mem[16'h1069] = 8'h01;
    mem[16'h106A] = 8'h81; // ADDN RSP 8
    mem[16'h106B] = 8'h06;
    mem[16'h106C] = 8'h08;
    mem[16'h106D] = 8'h00;
    mem[16'h106E] = 8'h00;
    mem[16'h106F] = 8'h00;
                          // .Lend8:
    mem[16'h1070] = 8'h40; // MOV RAX RBP
    mem[16'h1071] = 8'h00;
    mem[16'h1072] = 8'h05;
    mem[16'h1073] = 8'h85; // SUBN RAX 4
    mem[16'h1074] = 8'h00;
    mem[16'h1075] = 8'h04;
    mem[16'h1076] = 8'h00;
    mem[16'h1077] = 8'h00;
    mem[16'h1078] = 8'h00;
    mem[16'h1079] = 8'h85; // SUBN RSP 8
    mem[16'h107A] = 8'h06;
    mem[16'h107B] = 8'h08;
    mem[16'h107C] = 8'h00;
    mem[16'h107D] = 8'h00;
    mem[16'h107E] = 8'h00;
    mem[16'h107F] = 8'h04; // PUSH RAX
    mem[16'h1080] = 8'h00;
    mem[16'h1081] = 8'h85; // SUBN RSP 8
    mem[16'h1082] = 8'h06;
    mem[16'h1083] = 8'h08;
    mem[16'h1084] = 8'h00;
    mem[16'h1085] = 8'h00;
    mem[16'h1086] = 8'h00;
    mem[16'h1087] = 8'h05; // PUSHN 0
    mem[16'h1088] = 8'h00;
    mem[16'h1089] = 8'h00;
    mem[16'h108A] = 8'h00;
    mem[16'h108B] = 8'h00;
    mem[16'h108C] = 8'h00;
    mem[16'h108D] = 8'h08; // POP RDI
    mem[16'h108E] = 8'h01;
    mem[16'h108F] = 8'h81; // ADDN RSP 8
    mem[16'h1090] = 8'h06;
    mem[16'h1091] = 8'h08;
    mem[16'h1092] = 8'h00;
    mem[16'h1093] = 8'h00;
    mem[16'h1094] = 8'h00;
    mem[16'h1095] = 8'h08; // POP RAX
    mem[16'h1096] = 8'h00;
    mem[16'h1097] = 8'h81; // ADDN RSP 8
    mem[16'h1098] = 8'h06;
    mem[16'h1099] = 8'h08;
    mem[16'h109A] = 8'h00;
    mem[16'h109B] = 8'h00;
    mem[16'h109C] = 8'h00;
    mem[16'h109D] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h109E] = 8'h00;
    mem[16'h109F] = 8'h01;
    mem[16'h10A0] = 8'h85; // SUBN RSP 8
    mem[16'h10A1] = 8'h06;
    mem[16'h10A2] = 8'h08;
    mem[16'h10A3] = 8'h00;
    mem[16'h10A4] = 8'h00;
    mem[16'h10A5] = 8'h00;
    mem[16'h10A6] = 8'h04; // PUSH RDI
    mem[16'h10A7] = 8'h01;
    mem[16'h10A8] = 8'h81; // ADDN RSP 8
    mem[16'h10A9] = 8'h06;
    mem[16'h10AA] = 8'h08;
    mem[16'h10AB] = 8'h00;
    mem[16'h10AC] = 8'h00;
    mem[16'h10AD] = 8'h00;
                          // .Lbegin9:
    mem[16'h10AE] = 8'h40; // MOV RAX RBP
    mem[16'h10AF] = 8'h00;
    mem[16'h10B0] = 8'h05;
    mem[16'h10B1] = 8'h85; // SUBN RAX 4
    mem[16'h10B2] = 8'h00;
    mem[16'h10B3] = 8'h04;
    mem[16'h10B4] = 8'h00;
    mem[16'h10B5] = 8'h00;
    mem[16'h10B6] = 8'h00;
    mem[16'h10B7] = 8'h85; // SUBN RSP 8
    mem[16'h10B8] = 8'h06;
    mem[16'h10B9] = 8'h08;
    mem[16'h10BA] = 8'h00;
    mem[16'h10BB] = 8'h00;
    mem[16'h10BC] = 8'h00;
    mem[16'h10BD] = 8'h04; // PUSH RAX
    mem[16'h10BE] = 8'h00;
    mem[16'h10BF] = 8'h08; // POP RAX
    mem[16'h10C0] = 8'h00;
    mem[16'h10C1] = 8'h81; // ADDN RSP 8
    mem[16'h10C2] = 8'h06;
    mem[16'h10C3] = 8'h08;
    mem[16'h10C4] = 8'h00;
    mem[16'h10C5] = 8'h00;
    mem[16'h10C6] = 8'h00;
    mem[16'h10C7] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h10C8] = 8'h00;
    mem[16'h10C9] = 8'h00;
    mem[16'h10CA] = 8'h85; // SUBN RSP 8
    mem[16'h10CB] = 8'h06;
    mem[16'h10CC] = 8'h08;
    mem[16'h10CD] = 8'h00;
    mem[16'h10CE] = 8'h00;
    mem[16'h10CF] = 8'h00;
    mem[16'h10D0] = 8'h04; // PUSH RAX
    mem[16'h10D1] = 8'h00;
    mem[16'h10D2] = 8'h40; // MOV RAX RBP
    mem[16'h10D3] = 8'h00;
    mem[16'h10D4] = 8'h05;
    mem[16'h10D5] = 8'h85; // SUBN RAX 8
    mem[16'h10D6] = 8'h00;
    mem[16'h10D7] = 8'h08;
    mem[16'h10D8] = 8'h00;
    mem[16'h10D9] = 8'h00;
    mem[16'h10DA] = 8'h00;
    mem[16'h10DB] = 8'h85; // SUBN RSP 8
    mem[16'h10DC] = 8'h06;
    mem[16'h10DD] = 8'h08;
    mem[16'h10DE] = 8'h00;
    mem[16'h10DF] = 8'h00;
    mem[16'h10E0] = 8'h00;
    mem[16'h10E1] = 8'h04; // PUSH RAX
    mem[16'h10E2] = 8'h00;
    mem[16'h10E3] = 8'h08; // POP RAX
    mem[16'h10E4] = 8'h00;
    mem[16'h10E5] = 8'h81; // ADDN RSP 8
    mem[16'h10E6] = 8'h06;
    mem[16'h10E7] = 8'h08;
    mem[16'h10E8] = 8'h00;
    mem[16'h10E9] = 8'h00;
    mem[16'h10EA] = 8'h00;
    mem[16'h10EB] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h10EC] = 8'h00;
    mem[16'h10ED] = 8'h00;
    mem[16'h10EE] = 8'h85; // SUBN RSP 8
    mem[16'h10EF] = 8'h06;
    mem[16'h10F0] = 8'h08;
    mem[16'h10F1] = 8'h00;
    mem[16'h10F2] = 8'h00;
    mem[16'h10F3] = 8'h00;
    mem[16'h10F4] = 8'h04; // PUSH RAX
    mem[16'h10F5] = 8'h00;
    mem[16'h10F6] = 8'h08; // POP RDI
    mem[16'h10F7] = 8'h01;
    mem[16'h10F8] = 8'h81; // ADDN RSP 8
    mem[16'h10F9] = 8'h06;
    mem[16'h10FA] = 8'h08;
    mem[16'h10FB] = 8'h00;
    mem[16'h10FC] = 8'h00;
    mem[16'h10FD] = 8'h00;
    mem[16'h10FE] = 8'h08; // POP RAX
    mem[16'h10FF] = 8'h00;
    mem[16'h1100] = 8'h81; // ADDN RSP 8
    mem[16'h1101] = 8'h06;
    mem[16'h1102] = 8'h08;
    mem[16'h1103] = 8'h00;
    mem[16'h1104] = 8'h00;
    mem[16'h1105] = 8'h00;
    mem[16'h1106] = 8'h90; // CMP RAX RDI
    mem[16'h1107] = 8'h00;
    mem[16'h1108] = 8'h01;
    mem[16'h1109] = 8'h18; // SETL RAX
    mem[16'h110A] = 8'h00;
    mem[16'h110B] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h110C] = 8'h00;
    mem[16'h110D] = 8'h00;
    mem[16'h110E] = 8'h85; // SUBN RSP 8
    mem[16'h110F] = 8'h06;
    mem[16'h1110] = 8'h08;
    mem[16'h1111] = 8'h00;
    mem[16'h1112] = 8'h00;
    mem[16'h1113] = 8'h00;
    mem[16'h1114] = 8'h04; // PUSH RAX
    mem[16'h1115] = 8'h00;
    mem[16'h1116] = 8'h08; // POP RAX
    mem[16'h1117] = 8'h00;
    mem[16'h1118] = 8'h81; // ADDN RSP 8
    mem[16'h1119] = 8'h06;
    mem[16'h111A] = 8'h08;
    mem[16'h111B] = 8'h00;
    mem[16'h111C] = 8'h00;
    mem[16'h111D] = 8'h00;
    mem[16'h111E] = 8'h91; // CMPN RAX 0
    mem[16'h111F] = 8'h00;
    mem[16'h1120] = 8'h00;
    mem[16'h1121] = 8'h00;
    mem[16'h1122] = 8'h00;
    mem[16'h1123] = 8'h00;
    mem[16'h1124] = 8'h26; // JE .Lend9
    mem[16'h1125] = 8'hEB;
    mem[16'h1126] = 8'h15;
    mem[16'h1127] = 8'h00;
    mem[16'h1128] = 8'h00;
    mem[16'h1129] = 8'h00;
    mem[16'h112A] = 8'h00;
    mem[16'h112B] = 8'h00;
    mem[16'h112C] = 8'h00;
    mem[16'h112D] = 8'h40; // MOV RAX RBP
    mem[16'h112E] = 8'h00;
    mem[16'h112F] = 8'h05;
    mem[16'h1130] = 8'h85; // SUBN RAX 20
    mem[16'h1131] = 8'h00;
    mem[16'h1132] = 8'h14;
    mem[16'h1133] = 8'h00;
    mem[16'h1134] = 8'h00;
    mem[16'h1135] = 8'h00;
    mem[16'h1136] = 8'h85; // SUBN RSP 8
    mem[16'h1137] = 8'h06;
    mem[16'h1138] = 8'h08;
    mem[16'h1139] = 8'h00;
    mem[16'h113A] = 8'h00;
    mem[16'h113B] = 8'h00;
    mem[16'h113C] = 8'h04; // PUSH RAX
    mem[16'h113D] = 8'h00;
    mem[16'h113E] = 8'h85; // SUBN RSP 8
    mem[16'h113F] = 8'h06;
    mem[16'h1140] = 8'h08;
    mem[16'h1141] = 8'h00;
    mem[16'h1142] = 8'h00;
    mem[16'h1143] = 8'h00;
    mem[16'h1144] = 8'h05; // PUSHN 0
    mem[16'h1145] = 8'h00;
    mem[16'h1146] = 8'h00;
    mem[16'h1147] = 8'h00;
    mem[16'h1148] = 8'h00;
    mem[16'h1149] = 8'h00;
    mem[16'h114A] = 8'h08; // POP RDI
    mem[16'h114B] = 8'h01;
    mem[16'h114C] = 8'h81; // ADDN RSP 8
    mem[16'h114D] = 8'h06;
    mem[16'h114E] = 8'h08;
    mem[16'h114F] = 8'h00;
    mem[16'h1150] = 8'h00;
    mem[16'h1151] = 8'h00;
    mem[16'h1152] = 8'h08; // POP RAX
    mem[16'h1153] = 8'h00;
    mem[16'h1154] = 8'h81; // ADDN RSP 8
    mem[16'h1155] = 8'h06;
    mem[16'h1156] = 8'h08;
    mem[16'h1157] = 8'h00;
    mem[16'h1158] = 8'h00;
    mem[16'h1159] = 8'h00;
    mem[16'h115A] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h115B] = 8'h00;
    mem[16'h115C] = 8'h01;
    mem[16'h115D] = 8'h85; // SUBN RSP 8
    mem[16'h115E] = 8'h06;
    mem[16'h115F] = 8'h08;
    mem[16'h1160] = 8'h00;
    mem[16'h1161] = 8'h00;
    mem[16'h1162] = 8'h00;
    mem[16'h1163] = 8'h04; // PUSH RDI
    mem[16'h1164] = 8'h01;
    mem[16'h1165] = 8'h81; // ADDN RSP 8
    mem[16'h1166] = 8'h06;
    mem[16'h1167] = 8'h08;
    mem[16'h1168] = 8'h00;
    mem[16'h1169] = 8'h00;
    mem[16'h116A] = 8'h00;
                          // .Lbegin10:
    mem[16'h116B] = 8'h40; // MOV RAX RBP
    mem[16'h116C] = 8'h00;
    mem[16'h116D] = 8'h05;
    mem[16'h116E] = 8'h85; // SUBN RAX 20
    mem[16'h116F] = 8'h00;
    mem[16'h1170] = 8'h14;
    mem[16'h1171] = 8'h00;
    mem[16'h1172] = 8'h00;
    mem[16'h1173] = 8'h00;
    mem[16'h1174] = 8'h85; // SUBN RSP 8
    mem[16'h1175] = 8'h06;
    mem[16'h1176] = 8'h08;
    mem[16'h1177] = 8'h00;
    mem[16'h1178] = 8'h00;
    mem[16'h1179] = 8'h00;
    mem[16'h117A] = 8'h04; // PUSH RAX
    mem[16'h117B] = 8'h00;
    mem[16'h117C] = 8'h08; // POP RAX
    mem[16'h117D] = 8'h00;
    mem[16'h117E] = 8'h81; // ADDN RSP 8
    mem[16'h117F] = 8'h06;
    mem[16'h1180] = 8'h08;
    mem[16'h1181] = 8'h00;
    mem[16'h1182] = 8'h00;
    mem[16'h1183] = 8'h00;
    mem[16'h1184] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1185] = 8'h00;
    mem[16'h1186] = 8'h00;
    mem[16'h1187] = 8'h85; // SUBN RSP 8
    mem[16'h1188] = 8'h06;
    mem[16'h1189] = 8'h08;
    mem[16'h118A] = 8'h00;
    mem[16'h118B] = 8'h00;
    mem[16'h118C] = 8'h00;
    mem[16'h118D] = 8'h04; // PUSH RAX
    mem[16'h118E] = 8'h00;
    mem[16'h118F] = 8'h40; // MOV RAX RBP
    mem[16'h1190] = 8'h00;
    mem[16'h1191] = 8'h05;
    mem[16'h1192] = 8'h85; // SUBN RAX 24
    mem[16'h1193] = 8'h00;
    mem[16'h1194] = 8'h18;
    mem[16'h1195] = 8'h00;
    mem[16'h1196] = 8'h00;
    mem[16'h1197] = 8'h00;
    mem[16'h1198] = 8'h85; // SUBN RSP 8
    mem[16'h1199] = 8'h06;
    mem[16'h119A] = 8'h08;
    mem[16'h119B] = 8'h00;
    mem[16'h119C] = 8'h00;
    mem[16'h119D] = 8'h00;
    mem[16'h119E] = 8'h04; // PUSH RAX
    mem[16'h119F] = 8'h00;
    mem[16'h11A0] = 8'h08; // POP RAX
    mem[16'h11A1] = 8'h00;
    mem[16'h11A2] = 8'h81; // ADDN RSP 8
    mem[16'h11A3] = 8'h06;
    mem[16'h11A4] = 8'h08;
    mem[16'h11A5] = 8'h00;
    mem[16'h11A6] = 8'h00;
    mem[16'h11A7] = 8'h00;
    mem[16'h11A8] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h11A9] = 8'h00;
    mem[16'h11AA] = 8'h00;
    mem[16'h11AB] = 8'h85; // SUBN RSP 8
    mem[16'h11AC] = 8'h06;
    mem[16'h11AD] = 8'h08;
    mem[16'h11AE] = 8'h00;
    mem[16'h11AF] = 8'h00;
    mem[16'h11B0] = 8'h00;
    mem[16'h11B1] = 8'h04; // PUSH RAX
    mem[16'h11B2] = 8'h00;
    mem[16'h11B3] = 8'h08; // POP RDI
    mem[16'h11B4] = 8'h01;
    mem[16'h11B5] = 8'h81; // ADDN RSP 8
    mem[16'h11B6] = 8'h06;
    mem[16'h11B7] = 8'h08;
    mem[16'h11B8] = 8'h00;
    mem[16'h11B9] = 8'h00;
    mem[16'h11BA] = 8'h00;
    mem[16'h11BB] = 8'h08; // POP RAX
    mem[16'h11BC] = 8'h00;
    mem[16'h11BD] = 8'h81; // ADDN RSP 8
    mem[16'h11BE] = 8'h06;
    mem[16'h11BF] = 8'h08;
    mem[16'h11C0] = 8'h00;
    mem[16'h11C1] = 8'h00;
    mem[16'h11C2] = 8'h00;
    mem[16'h11C3] = 8'h90; // CMP RAX RDI
    mem[16'h11C4] = 8'h00;
    mem[16'h11C5] = 8'h01;
    mem[16'h11C6] = 8'h18; // SETL RAX
    mem[16'h11C7] = 8'h00;
    mem[16'h11C8] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h11C9] = 8'h00;
    mem[16'h11CA] = 8'h00;
    mem[16'h11CB] = 8'h85; // SUBN RSP 8
    mem[16'h11CC] = 8'h06;
    mem[16'h11CD] = 8'h08;
    mem[16'h11CE] = 8'h00;
    mem[16'h11CF] = 8'h00;
    mem[16'h11D0] = 8'h00;
    mem[16'h11D1] = 8'h04; // PUSH RAX
    mem[16'h11D2] = 8'h00;
    mem[16'h11D3] = 8'h08; // POP RAX
    mem[16'h11D4] = 8'h00;
    mem[16'h11D5] = 8'h81; // ADDN RSP 8
    mem[16'h11D6] = 8'h06;
    mem[16'h11D7] = 8'h08;
    mem[16'h11D8] = 8'h00;
    mem[16'h11D9] = 8'h00;
    mem[16'h11DA] = 8'h00;
    mem[16'h11DB] = 8'h91; // CMPN RAX 0
    mem[16'h11DC] = 8'h00;
    mem[16'h11DD] = 8'h00;
    mem[16'h11DE] = 8'h00;
    mem[16'h11DF] = 8'h00;
    mem[16'h11E0] = 8'h00;
    mem[16'h11E1] = 8'h26; // JE .Lend10
    mem[16'h11E2] = 8'h6B;
    mem[16'h11E3] = 8'h14;
    mem[16'h11E4] = 8'h00;
    mem[16'h11E5] = 8'h00;
    mem[16'h11E6] = 8'h00;
    mem[16'h11E7] = 8'h00;
    mem[16'h11E8] = 8'h00;
    mem[16'h11E9] = 8'h00;
    mem[16'h11EA] = 8'h85; // SUBN RSP 8
    mem[16'h11EB] = 8'h06;
    mem[16'h11EC] = 8'h08;
    mem[16'h11ED] = 8'h00;
    mem[16'h11EE] = 8'h00;
    mem[16'h11EF] = 8'h00;
    mem[16'h11F0] = 8'h06; // PUSHA pos
    mem[16'h11F1] = 8'h09;
    mem[16'h11F2] = 8'h00;
    mem[16'h11F3] = 8'h00;
    mem[16'h11F4] = 8'h00;
    mem[16'h11F5] = 8'h00;
    mem[16'h11F6] = 8'h00;
    mem[16'h11F7] = 8'h00;
    mem[16'h11F8] = 8'h00;
    mem[16'h11F9] = 8'h40; // MOV RAX RBP
    mem[16'h11FA] = 8'h00;
    mem[16'h11FB] = 8'h05;
    mem[16'h11FC] = 8'h85; // SUBN RAX 20
    mem[16'h11FD] = 8'h00;
    mem[16'h11FE] = 8'h14;
    mem[16'h11FF] = 8'h00;
    mem[16'h1200] = 8'h00;
    mem[16'h1201] = 8'h00;
    mem[16'h1202] = 8'h85; // SUBN RSP 8
    mem[16'h1203] = 8'h06;
    mem[16'h1204] = 8'h08;
    mem[16'h1205] = 8'h00;
    mem[16'h1206] = 8'h00;
    mem[16'h1207] = 8'h00;
    mem[16'h1208] = 8'h04; // PUSH RAX
    mem[16'h1209] = 8'h00;
    mem[16'h120A] = 8'h08; // POP RAX
    mem[16'h120B] = 8'h00;
    mem[16'h120C] = 8'h81; // ADDN RSP 8
    mem[16'h120D] = 8'h06;
    mem[16'h120E] = 8'h08;
    mem[16'h120F] = 8'h00;
    mem[16'h1210] = 8'h00;
    mem[16'h1211] = 8'h00;
    mem[16'h1212] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1213] = 8'h00;
    mem[16'h1214] = 8'h00;
    mem[16'h1215] = 8'h85; // SUBN RSP 8
    mem[16'h1216] = 8'h06;
    mem[16'h1217] = 8'h08;
    mem[16'h1218] = 8'h00;
    mem[16'h1219] = 8'h00;
    mem[16'h121A] = 8'h00;
    mem[16'h121B] = 8'h04; // PUSH RAX
    mem[16'h121C] = 8'h00;
    mem[16'h121D] = 8'h08; // POP RDI
    mem[16'h121E] = 8'h01;
    mem[16'h121F] = 8'h81; // ADDN RSP 8
    mem[16'h1220] = 8'h06;
    mem[16'h1221] = 8'h08;
    mem[16'h1222] = 8'h00;
    mem[16'h1223] = 8'h00;
    mem[16'h1224] = 8'h00;
    mem[16'h1225] = 8'h08; // POP RAX
    mem[16'h1226] = 8'h00;
    mem[16'h1227] = 8'h81; // ADDN RSP 8
    mem[16'h1228] = 8'h06;
    mem[16'h1229] = 8'h08;
    mem[16'h122A] = 8'h00;
    mem[16'h122B] = 8'h00;
    mem[16'h122C] = 8'h00;
    mem[16'h122D] = 8'h89; // MULN RDI 8
    mem[16'h122E] = 8'h01;
    mem[16'h122F] = 8'h08;
    mem[16'h1230] = 8'h00;
    mem[16'h1231] = 8'h00;
    mem[16'h1232] = 8'h00;
    mem[16'h1233] = 8'h80; // ADD RAX RDI
    mem[16'h1234] = 8'h00;
    mem[16'h1235] = 8'h01;
    mem[16'h1236] = 8'h85; // SUBN RSP 8
    mem[16'h1237] = 8'h06;
    mem[16'h1238] = 8'h08;
    mem[16'h1239] = 8'h00;
    mem[16'h123A] = 8'h00;
    mem[16'h123B] = 8'h00;
    mem[16'h123C] = 8'h04; // PUSH RAX
    mem[16'h123D] = 8'h00;
    mem[16'h123E] = 8'h85; // SUBN RSP 8
    mem[16'h123F] = 8'h06;
    mem[16'h1240] = 8'h08;
    mem[16'h1241] = 8'h00;
    mem[16'h1242] = 8'h00;
    mem[16'h1243] = 8'h00;
    mem[16'h1244] = 8'h05; // PUSHN 0
    mem[16'h1245] = 8'h00;
    mem[16'h1246] = 8'h00;
    mem[16'h1247] = 8'h00;
    mem[16'h1248] = 8'h00;
    mem[16'h1249] = 8'h00;
    mem[16'h124A] = 8'h08; // POP RDI
    mem[16'h124B] = 8'h01;
    mem[16'h124C] = 8'h81; // ADDN RSP 8
    mem[16'h124D] = 8'h06;
    mem[16'h124E] = 8'h08;
    mem[16'h124F] = 8'h00;
    mem[16'h1250] = 8'h00;
    mem[16'h1251] = 8'h00;
    mem[16'h1252] = 8'h08; // POP RAX
    mem[16'h1253] = 8'h00;
    mem[16'h1254] = 8'h81; // ADDN RSP 8
    mem[16'h1255] = 8'h06;
    mem[16'h1256] = 8'h08;
    mem[16'h1257] = 8'h00;
    mem[16'h1258] = 8'h00;
    mem[16'h1259] = 8'h00;
    mem[16'h125A] = 8'h89; // MULN RDI 4
    mem[16'h125B] = 8'h01;
    mem[16'h125C] = 8'h04;
    mem[16'h125D] = 8'h00;
    mem[16'h125E] = 8'h00;
    mem[16'h125F] = 8'h00;
    mem[16'h1260] = 8'h80; // ADD RAX RDI
    mem[16'h1261] = 8'h00;
    mem[16'h1262] = 8'h01;
    mem[16'h1263] = 8'h85; // SUBN RSP 8
    mem[16'h1264] = 8'h06;
    mem[16'h1265] = 8'h08;
    mem[16'h1266] = 8'h00;
    mem[16'h1267] = 8'h00;
    mem[16'h1268] = 8'h00;
    mem[16'h1269] = 8'h04; // PUSH RAX
    mem[16'h126A] = 8'h00;
    mem[16'h126B] = 8'h08; // POP RAX
    mem[16'h126C] = 8'h00;
    mem[16'h126D] = 8'h81; // ADDN RSP 8
    mem[16'h126E] = 8'h06;
    mem[16'h126F] = 8'h08;
    mem[16'h1270] = 8'h00;
    mem[16'h1271] = 8'h00;
    mem[16'h1272] = 8'h00;
    mem[16'h1273] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1274] = 8'h00;
    mem[16'h1275] = 8'h00;
    mem[16'h1276] = 8'h85; // SUBN RSP 8
    mem[16'h1277] = 8'h06;
    mem[16'h1278] = 8'h08;
    mem[16'h1279] = 8'h00;
    mem[16'h127A] = 8'h00;
    mem[16'h127B] = 8'h00;
    mem[16'h127C] = 8'h04; // PUSH RAX
    mem[16'h127D] = 8'h00;
    mem[16'h127E] = 8'h40; // MOV RAX RBP
    mem[16'h127F] = 8'h00;
    mem[16'h1280] = 8'h05;
    mem[16'h1281] = 8'h85; // SUBN RAX 16
    mem[16'h1282] = 8'h00;
    mem[16'h1283] = 8'h10;
    mem[16'h1284] = 8'h00;
    mem[16'h1285] = 8'h00;
    mem[16'h1286] = 8'h00;
    mem[16'h1287] = 8'h85; // SUBN RSP 8
    mem[16'h1288] = 8'h06;
    mem[16'h1289] = 8'h08;
    mem[16'h128A] = 8'h00;
    mem[16'h128B] = 8'h00;
    mem[16'h128C] = 8'h00;
    mem[16'h128D] = 8'h04; // PUSH RAX
    mem[16'h128E] = 8'h00;
    mem[16'h128F] = 8'h08; // POP RAX
    mem[16'h1290] = 8'h00;
    mem[16'h1291] = 8'h81; // ADDN RSP 8
    mem[16'h1292] = 8'h06;
    mem[16'h1293] = 8'h08;
    mem[16'h1294] = 8'h00;
    mem[16'h1295] = 8'h00;
    mem[16'h1296] = 8'h00;
    mem[16'h1297] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1298] = 8'h00;
    mem[16'h1299] = 8'h00;
    mem[16'h129A] = 8'h85; // SUBN RSP 8
    mem[16'h129B] = 8'h06;
    mem[16'h129C] = 8'h08;
    mem[16'h129D] = 8'h00;
    mem[16'h129E] = 8'h00;
    mem[16'h129F] = 8'h00;
    mem[16'h12A0] = 8'h04; // PUSH RAX
    mem[16'h12A1] = 8'h00;
    mem[16'h12A2] = 8'h08; // POP RDI
    mem[16'h12A3] = 8'h01;
    mem[16'h12A4] = 8'h81; // ADDN RSP 8
    mem[16'h12A5] = 8'h06;
    mem[16'h12A6] = 8'h08;
    mem[16'h12A7] = 8'h00;
    mem[16'h12A8] = 8'h00;
    mem[16'h12A9] = 8'h00;
    mem[16'h12AA] = 8'h08; // POP RAX
    mem[16'h12AB] = 8'h00;
    mem[16'h12AC] = 8'h81; // ADDN RSP 8
    mem[16'h12AD] = 8'h06;
    mem[16'h12AE] = 8'h08;
    mem[16'h12AF] = 8'h00;
    mem[16'h12B0] = 8'h00;
    mem[16'h12B1] = 8'h00;
    mem[16'h12B2] = 8'h90; // CMP RAX RDI
    mem[16'h12B3] = 8'h00;
    mem[16'h12B4] = 8'h01;
    mem[16'h12B5] = 8'h10; // SETE RAX
    mem[16'h12B6] = 8'h00;
    mem[16'h12B7] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h12B8] = 8'h00;
    mem[16'h12B9] = 8'h00;
    mem[16'h12BA] = 8'h85; // SUBN RSP 8
    mem[16'h12BB] = 8'h06;
    mem[16'h12BC] = 8'h08;
    mem[16'h12BD] = 8'h00;
    mem[16'h12BE] = 8'h00;
    mem[16'h12BF] = 8'h00;
    mem[16'h12C0] = 8'h04; // PUSH RAX
    mem[16'h12C1] = 8'h00;
    mem[16'h12C2] = 8'h08; // POP RAX
    mem[16'h12C3] = 8'h00;
    mem[16'h12C4] = 8'h81; // ADDN RSP 8
    mem[16'h12C5] = 8'h06;
    mem[16'h12C6] = 8'h08;
    mem[16'h12C7] = 8'h00;
    mem[16'h12C8] = 8'h00;
    mem[16'h12C9] = 8'h00;
    mem[16'h12CA] = 8'h91; // CMPN RAX 0
    mem[16'h12CB] = 8'h00;
    mem[16'h12CC] = 8'h00;
    mem[16'h12CD] = 8'h00;
    mem[16'h12CE] = 8'h00;
    mem[16'h12CF] = 8'h00;
    mem[16'h12D0] = 8'h26; // JE .Lend11
    mem[16'h12D1] = 8'hE5;
    mem[16'h12D2] = 8'h13;
    mem[16'h12D3] = 8'h00;
    mem[16'h12D4] = 8'h00;
    mem[16'h12D5] = 8'h00;
    mem[16'h12D6] = 8'h00;
    mem[16'h12D7] = 8'h00;
    mem[16'h12D8] = 8'h00;
    mem[16'h12D9] = 8'h85; // SUBN RSP 8
    mem[16'h12DA] = 8'h06;
    mem[16'h12DB] = 8'h08;
    mem[16'h12DC] = 8'h00;
    mem[16'h12DD] = 8'h00;
    mem[16'h12DE] = 8'h00;
    mem[16'h12DF] = 8'h06; // PUSHA pos
    mem[16'h12E0] = 8'h09;
    mem[16'h12E1] = 8'h00;
    mem[16'h12E2] = 8'h00;
    mem[16'h12E3] = 8'h00;
    mem[16'h12E4] = 8'h00;
    mem[16'h12E5] = 8'h00;
    mem[16'h12E6] = 8'h00;
    mem[16'h12E7] = 8'h00;
    mem[16'h12E8] = 8'h40; // MOV RAX RBP
    mem[16'h12E9] = 8'h00;
    mem[16'h12EA] = 8'h05;
    mem[16'h12EB] = 8'h85; // SUBN RAX 20
    mem[16'h12EC] = 8'h00;
    mem[16'h12ED] = 8'h14;
    mem[16'h12EE] = 8'h00;
    mem[16'h12EF] = 8'h00;
    mem[16'h12F0] = 8'h00;
    mem[16'h12F1] = 8'h85; // SUBN RSP 8
    mem[16'h12F2] = 8'h06;
    mem[16'h12F3] = 8'h08;
    mem[16'h12F4] = 8'h00;
    mem[16'h12F5] = 8'h00;
    mem[16'h12F6] = 8'h00;
    mem[16'h12F7] = 8'h04; // PUSH RAX
    mem[16'h12F8] = 8'h00;
    mem[16'h12F9] = 8'h08; // POP RAX
    mem[16'h12FA] = 8'h00;
    mem[16'h12FB] = 8'h81; // ADDN RSP 8
    mem[16'h12FC] = 8'h06;
    mem[16'h12FD] = 8'h08;
    mem[16'h12FE] = 8'h00;
    mem[16'h12FF] = 8'h00;
    mem[16'h1300] = 8'h00;
    mem[16'h1301] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1302] = 8'h00;
    mem[16'h1303] = 8'h00;
    mem[16'h1304] = 8'h85; // SUBN RSP 8
    mem[16'h1305] = 8'h06;
    mem[16'h1306] = 8'h08;
    mem[16'h1307] = 8'h00;
    mem[16'h1308] = 8'h00;
    mem[16'h1309] = 8'h00;
    mem[16'h130A] = 8'h04; // PUSH RAX
    mem[16'h130B] = 8'h00;
    mem[16'h130C] = 8'h08; // POP RDI
    mem[16'h130D] = 8'h01;
    mem[16'h130E] = 8'h81; // ADDN RSP 8
    mem[16'h130F] = 8'h06;
    mem[16'h1310] = 8'h08;
    mem[16'h1311] = 8'h00;
    mem[16'h1312] = 8'h00;
    mem[16'h1313] = 8'h00;
    mem[16'h1314] = 8'h08; // POP RAX
    mem[16'h1315] = 8'h00;
    mem[16'h1316] = 8'h81; // ADDN RSP 8
    mem[16'h1317] = 8'h06;
    mem[16'h1318] = 8'h08;
    mem[16'h1319] = 8'h00;
    mem[16'h131A] = 8'h00;
    mem[16'h131B] = 8'h00;
    mem[16'h131C] = 8'h89; // MULN RDI 8
    mem[16'h131D] = 8'h01;
    mem[16'h131E] = 8'h08;
    mem[16'h131F] = 8'h00;
    mem[16'h1320] = 8'h00;
    mem[16'h1321] = 8'h00;
    mem[16'h1322] = 8'h80; // ADD RAX RDI
    mem[16'h1323] = 8'h00;
    mem[16'h1324] = 8'h01;
    mem[16'h1325] = 8'h85; // SUBN RSP 8
    mem[16'h1326] = 8'h06;
    mem[16'h1327] = 8'h08;
    mem[16'h1328] = 8'h00;
    mem[16'h1329] = 8'h00;
    mem[16'h132A] = 8'h00;
    mem[16'h132B] = 8'h04; // PUSH RAX
    mem[16'h132C] = 8'h00;
    mem[16'h132D] = 8'h85; // SUBN RSP 8
    mem[16'h132E] = 8'h06;
    mem[16'h132F] = 8'h08;
    mem[16'h1330] = 8'h00;
    mem[16'h1331] = 8'h00;
    mem[16'h1332] = 8'h00;
    mem[16'h1333] = 8'h05; // PUSHN 1
    mem[16'h1334] = 8'h00;
    mem[16'h1335] = 8'h01;
    mem[16'h1336] = 8'h00;
    mem[16'h1337] = 8'h00;
    mem[16'h1338] = 8'h00;
    mem[16'h1339] = 8'h08; // POP RDI
    mem[16'h133A] = 8'h01;
    mem[16'h133B] = 8'h81; // ADDN RSP 8
    mem[16'h133C] = 8'h06;
    mem[16'h133D] = 8'h08;
    mem[16'h133E] = 8'h00;
    mem[16'h133F] = 8'h00;
    mem[16'h1340] = 8'h00;
    mem[16'h1341] = 8'h08; // POP RAX
    mem[16'h1342] = 8'h00;
    mem[16'h1343] = 8'h81; // ADDN RSP 8
    mem[16'h1344] = 8'h06;
    mem[16'h1345] = 8'h08;
    mem[16'h1346] = 8'h00;
    mem[16'h1347] = 8'h00;
    mem[16'h1348] = 8'h00;
    mem[16'h1349] = 8'h89; // MULN RDI 4
    mem[16'h134A] = 8'h01;
    mem[16'h134B] = 8'h04;
    mem[16'h134C] = 8'h00;
    mem[16'h134D] = 8'h00;
    mem[16'h134E] = 8'h00;
    mem[16'h134F] = 8'h80; // ADD RAX RDI
    mem[16'h1350] = 8'h00;
    mem[16'h1351] = 8'h01;
    mem[16'h1352] = 8'h85; // SUBN RSP 8
    mem[16'h1353] = 8'h06;
    mem[16'h1354] = 8'h08;
    mem[16'h1355] = 8'h00;
    mem[16'h1356] = 8'h00;
    mem[16'h1357] = 8'h00;
    mem[16'h1358] = 8'h04; // PUSH RAX
    mem[16'h1359] = 8'h00;
    mem[16'h135A] = 8'h08; // POP RAX
    mem[16'h135B] = 8'h00;
    mem[16'h135C] = 8'h81; // ADDN RSP 8
    mem[16'h135D] = 8'h06;
    mem[16'h135E] = 8'h08;
    mem[16'h135F] = 8'h00;
    mem[16'h1360] = 8'h00;
    mem[16'h1361] = 8'h00;
    mem[16'h1362] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1363] = 8'h00;
    mem[16'h1364] = 8'h00;
    mem[16'h1365] = 8'h85; // SUBN RSP 8
    mem[16'h1366] = 8'h06;
    mem[16'h1367] = 8'h08;
    mem[16'h1368] = 8'h00;
    mem[16'h1369] = 8'h00;
    mem[16'h136A] = 8'h00;
    mem[16'h136B] = 8'h04; // PUSH RAX
    mem[16'h136C] = 8'h00;
    mem[16'h136D] = 8'h40; // MOV RAX RBP
    mem[16'h136E] = 8'h00;
    mem[16'h136F] = 8'h05;
    mem[16'h1370] = 8'h85; // SUBN RAX 12
    mem[16'h1371] = 8'h00;
    mem[16'h1372] = 8'h0C;
    mem[16'h1373] = 8'h00;
    mem[16'h1374] = 8'h00;
    mem[16'h1375] = 8'h00;
    mem[16'h1376] = 8'h85; // SUBN RSP 8
    mem[16'h1377] = 8'h06;
    mem[16'h1378] = 8'h08;
    mem[16'h1379] = 8'h00;
    mem[16'h137A] = 8'h00;
    mem[16'h137B] = 8'h00;
    mem[16'h137C] = 8'h04; // PUSH RAX
    mem[16'h137D] = 8'h00;
    mem[16'h137E] = 8'h08; // POP RAX
    mem[16'h137F] = 8'h00;
    mem[16'h1380] = 8'h81; // ADDN RSP 8
    mem[16'h1381] = 8'h06;
    mem[16'h1382] = 8'h08;
    mem[16'h1383] = 8'h00;
    mem[16'h1384] = 8'h00;
    mem[16'h1385] = 8'h00;
    mem[16'h1386] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1387] = 8'h00;
    mem[16'h1388] = 8'h00;
    mem[16'h1389] = 8'h85; // SUBN RSP 8
    mem[16'h138A] = 8'h06;
    mem[16'h138B] = 8'h08;
    mem[16'h138C] = 8'h00;
    mem[16'h138D] = 8'h00;
    mem[16'h138E] = 8'h00;
    mem[16'h138F] = 8'h04; // PUSH RAX
    mem[16'h1390] = 8'h00;
    mem[16'h1391] = 8'h08; // POP RDI
    mem[16'h1392] = 8'h01;
    mem[16'h1393] = 8'h81; // ADDN RSP 8
    mem[16'h1394] = 8'h06;
    mem[16'h1395] = 8'h08;
    mem[16'h1396] = 8'h00;
    mem[16'h1397] = 8'h00;
    mem[16'h1398] = 8'h00;
    mem[16'h1399] = 8'h08; // POP RAX
    mem[16'h139A] = 8'h00;
    mem[16'h139B] = 8'h81; // ADDN RSP 8
    mem[16'h139C] = 8'h06;
    mem[16'h139D] = 8'h08;
    mem[16'h139E] = 8'h00;
    mem[16'h139F] = 8'h00;
    mem[16'h13A0] = 8'h00;
    mem[16'h13A1] = 8'h90; // CMP RAX RDI
    mem[16'h13A2] = 8'h00;
    mem[16'h13A3] = 8'h01;
    mem[16'h13A4] = 8'h10; // SETE RAX
    mem[16'h13A5] = 8'h00;
    mem[16'h13A6] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h13A7] = 8'h00;
    mem[16'h13A8] = 8'h00;
    mem[16'h13A9] = 8'h85; // SUBN RSP 8
    mem[16'h13AA] = 8'h06;
    mem[16'h13AB] = 8'h08;
    mem[16'h13AC] = 8'h00;
    mem[16'h13AD] = 8'h00;
    mem[16'h13AE] = 8'h00;
    mem[16'h13AF] = 8'h04; // PUSH RAX
    mem[16'h13B0] = 8'h00;
    mem[16'h13B1] = 8'h08; // POP RAX
    mem[16'h13B2] = 8'h00;
    mem[16'h13B3] = 8'h81; // ADDN RSP 8
    mem[16'h13B4] = 8'h06;
    mem[16'h13B5] = 8'h08;
    mem[16'h13B6] = 8'h00;
    mem[16'h13B7] = 8'h00;
    mem[16'h13B8] = 8'h00;
    mem[16'h13B9] = 8'h91; // CMPN RAX 0
    mem[16'h13BA] = 8'h00;
    mem[16'h13BB] = 8'h00;
    mem[16'h13BC] = 8'h00;
    mem[16'h13BD] = 8'h00;
    mem[16'h13BE] = 8'h00;
    mem[16'h13BF] = 8'h26; // JE .Lend12
    mem[16'h13C0] = 8'hE5;
    mem[16'h13C1] = 8'h13;
    mem[16'h13C2] = 8'h00;
    mem[16'h13C3] = 8'h00;
    mem[16'h13C4] = 8'h00;
    mem[16'h13C5] = 8'h00;
    mem[16'h13C6] = 8'h00;
    mem[16'h13C7] = 8'h00;
    mem[16'h13C8] = 8'h85; // SUBN RSP 8
    mem[16'h13C9] = 8'h06;
    mem[16'h13CA] = 8'h08;
    mem[16'h13CB] = 8'h00;
    mem[16'h13CC] = 8'h00;
    mem[16'h13CD] = 8'h00;
    mem[16'h13CE] = 8'h05; // PUSHN 0
    mem[16'h13CF] = 8'h00;
    mem[16'h13D0] = 8'h00;
    mem[16'h13D1] = 8'h00;
    mem[16'h13D2] = 8'h00;
    mem[16'h13D3] = 8'h00;
    mem[16'h13D4] = 8'h08; // POP RAX
    mem[16'h13D5] = 8'h00;
    mem[16'h13D6] = 8'h81; // ADDN RSP 8
    mem[16'h13D7] = 8'h06;
    mem[16'h13D8] = 8'h08;
    mem[16'h13D9] = 8'h00;
    mem[16'h13DA] = 8'h00;
    mem[16'h13DB] = 8'h00;
    mem[16'h13DC] = 8'h22; // JMP .Lreturn.check
    mem[16'h13DD] = 8'h08;
    mem[16'h13DE] = 8'h16;
    mem[16'h13DF] = 8'h00;
    mem[16'h13E0] = 8'h00;
    mem[16'h13E1] = 8'h00;
    mem[16'h13E2] = 8'h00;
    mem[16'h13E3] = 8'h00;
    mem[16'h13E4] = 8'h00;
                          // .Lend12:
                          // .Lend11:
    mem[16'h13E5] = 8'h40; // MOV RAX RBP
    mem[16'h13E6] = 8'h00;
    mem[16'h13E7] = 8'h05;
    mem[16'h13E8] = 8'h85; // SUBN RAX 20
    mem[16'h13E9] = 8'h00;
    mem[16'h13EA] = 8'h14;
    mem[16'h13EB] = 8'h00;
    mem[16'h13EC] = 8'h00;
    mem[16'h13ED] = 8'h00;
    mem[16'h13EE] = 8'h85; // SUBN RSP 8
    mem[16'h13EF] = 8'h06;
    mem[16'h13F0] = 8'h08;
    mem[16'h13F1] = 8'h00;
    mem[16'h13F2] = 8'h00;
    mem[16'h13F3] = 8'h00;
    mem[16'h13F4] = 8'h04; // PUSH RAX
    mem[16'h13F5] = 8'h00;
    mem[16'h13F6] = 8'h40; // MOV RAX RBP
    mem[16'h13F7] = 8'h00;
    mem[16'h13F8] = 8'h05;
    mem[16'h13F9] = 8'h85; // SUBN RAX 20
    mem[16'h13FA] = 8'h00;
    mem[16'h13FB] = 8'h14;
    mem[16'h13FC] = 8'h00;
    mem[16'h13FD] = 8'h00;
    mem[16'h13FE] = 8'h00;
    mem[16'h13FF] = 8'h85; // SUBN RSP 8
    mem[16'h1400] = 8'h06;
    mem[16'h1401] = 8'h08;
    mem[16'h1402] = 8'h00;
    mem[16'h1403] = 8'h00;
    mem[16'h1404] = 8'h00;
    mem[16'h1405] = 8'h04; // PUSH RAX
    mem[16'h1406] = 8'h00;
    mem[16'h1407] = 8'h08; // POP RAX
    mem[16'h1408] = 8'h00;
    mem[16'h1409] = 8'h81; // ADDN RSP 8
    mem[16'h140A] = 8'h06;
    mem[16'h140B] = 8'h08;
    mem[16'h140C] = 8'h00;
    mem[16'h140D] = 8'h00;
    mem[16'h140E] = 8'h00;
    mem[16'h140F] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1410] = 8'h00;
    mem[16'h1411] = 8'h00;
    mem[16'h1412] = 8'h85; // SUBN RSP 8
    mem[16'h1413] = 8'h06;
    mem[16'h1414] = 8'h08;
    mem[16'h1415] = 8'h00;
    mem[16'h1416] = 8'h00;
    mem[16'h1417] = 8'h00;
    mem[16'h1418] = 8'h04; // PUSH RAX
    mem[16'h1419] = 8'h00;
    mem[16'h141A] = 8'h85; // SUBN RSP 8
    mem[16'h141B] = 8'h06;
    mem[16'h141C] = 8'h08;
    mem[16'h141D] = 8'h00;
    mem[16'h141E] = 8'h00;
    mem[16'h141F] = 8'h00;
    mem[16'h1420] = 8'h05; // PUSHN 1
    mem[16'h1421] = 8'h00;
    mem[16'h1422] = 8'h01;
    mem[16'h1423] = 8'h00;
    mem[16'h1424] = 8'h00;
    mem[16'h1425] = 8'h00;
    mem[16'h1426] = 8'h08; // POP RDI
    mem[16'h1427] = 8'h01;
    mem[16'h1428] = 8'h81; // ADDN RSP 8
    mem[16'h1429] = 8'h06;
    mem[16'h142A] = 8'h08;
    mem[16'h142B] = 8'h00;
    mem[16'h142C] = 8'h00;
    mem[16'h142D] = 8'h00;
    mem[16'h142E] = 8'h08; // POP RAX
    mem[16'h142F] = 8'h00;
    mem[16'h1430] = 8'h81; // ADDN RSP 8
    mem[16'h1431] = 8'h06;
    mem[16'h1432] = 8'h08;
    mem[16'h1433] = 8'h00;
    mem[16'h1434] = 8'h00;
    mem[16'h1435] = 8'h00;
    mem[16'h1436] = 8'h80; // ADD RAX RDI
    mem[16'h1437] = 8'h00;
    mem[16'h1438] = 8'h01;
    mem[16'h1439] = 8'h85; // SUBN RSP 8
    mem[16'h143A] = 8'h06;
    mem[16'h143B] = 8'h08;
    mem[16'h143C] = 8'h00;
    mem[16'h143D] = 8'h00;
    mem[16'h143E] = 8'h00;
    mem[16'h143F] = 8'h04; // PUSH RAX
    mem[16'h1440] = 8'h00;
    mem[16'h1441] = 8'h08; // POP RDI
    mem[16'h1442] = 8'h01;
    mem[16'h1443] = 8'h81; // ADDN RSP 8
    mem[16'h1444] = 8'h06;
    mem[16'h1445] = 8'h08;
    mem[16'h1446] = 8'h00;
    mem[16'h1447] = 8'h00;
    mem[16'h1448] = 8'h00;
    mem[16'h1449] = 8'h08; // POP RAX
    mem[16'h144A] = 8'h00;
    mem[16'h144B] = 8'h81; // ADDN RSP 8
    mem[16'h144C] = 8'h06;
    mem[16'h144D] = 8'h08;
    mem[16'h144E] = 8'h00;
    mem[16'h144F] = 8'h00;
    mem[16'h1450] = 8'h00;
    mem[16'h1451] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h1452] = 8'h00;
    mem[16'h1453] = 8'h01;
    mem[16'h1454] = 8'h85; // SUBN RSP 8
    mem[16'h1455] = 8'h06;
    mem[16'h1456] = 8'h08;
    mem[16'h1457] = 8'h00;
    mem[16'h1458] = 8'h00;
    mem[16'h1459] = 8'h00;
    mem[16'h145A] = 8'h04; // PUSH RDI
    mem[16'h145B] = 8'h01;
    mem[16'h145C] = 8'h81; // ADDN RSP 8
    mem[16'h145D] = 8'h06;
    mem[16'h145E] = 8'h08;
    mem[16'h145F] = 8'h00;
    mem[16'h1460] = 8'h00;
    mem[16'h1461] = 8'h00;
    mem[16'h1462] = 8'h22; // JMP .Lbegin10
    mem[16'h1463] = 8'h6B;
    mem[16'h1464] = 8'h11;
    mem[16'h1465] = 8'h00;
    mem[16'h1466] = 8'h00;
    mem[16'h1467] = 8'h00;
    mem[16'h1468] = 8'h00;
    mem[16'h1469] = 8'h00;
    mem[16'h146A] = 8'h00;
                          // .Lend10:
    mem[16'h146B] = 8'h40; // MOV RAX RBP
    mem[16'h146C] = 8'h00;
    mem[16'h146D] = 8'h05;
    mem[16'h146E] = 8'h85; // SUBN RAX 16
    mem[16'h146F] = 8'h00;
    mem[16'h1470] = 8'h10;
    mem[16'h1471] = 8'h00;
    mem[16'h1472] = 8'h00;
    mem[16'h1473] = 8'h00;
    mem[16'h1474] = 8'h85; // SUBN RSP 8
    mem[16'h1475] = 8'h06;
    mem[16'h1476] = 8'h08;
    mem[16'h1477] = 8'h00;
    mem[16'h1478] = 8'h00;
    mem[16'h1479] = 8'h00;
    mem[16'h147A] = 8'h04; // PUSH RAX
    mem[16'h147B] = 8'h00;
    mem[16'h147C] = 8'h40; // MOV RAX RBP
    mem[16'h147D] = 8'h00;
    mem[16'h147E] = 8'h05;
    mem[16'h147F] = 8'h85; // SUBN RAX 16
    mem[16'h1480] = 8'h00;
    mem[16'h1481] = 8'h10;
    mem[16'h1482] = 8'h00;
    mem[16'h1483] = 8'h00;
    mem[16'h1484] = 8'h00;
    mem[16'h1485] = 8'h85; // SUBN RSP 8
    mem[16'h1486] = 8'h06;
    mem[16'h1487] = 8'h08;
    mem[16'h1488] = 8'h00;
    mem[16'h1489] = 8'h00;
    mem[16'h148A] = 8'h00;
    mem[16'h148B] = 8'h04; // PUSH RAX
    mem[16'h148C] = 8'h00;
    mem[16'h148D] = 8'h08; // POP RAX
    mem[16'h148E] = 8'h00;
    mem[16'h148F] = 8'h81; // ADDN RSP 8
    mem[16'h1490] = 8'h06;
    mem[16'h1491] = 8'h08;
    mem[16'h1492] = 8'h00;
    mem[16'h1493] = 8'h00;
    mem[16'h1494] = 8'h00;
    mem[16'h1495] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1496] = 8'h00;
    mem[16'h1497] = 8'h00;
    mem[16'h1498] = 8'h85; // SUBN RSP 8
    mem[16'h1499] = 8'h06;
    mem[16'h149A] = 8'h08;
    mem[16'h149B] = 8'h00;
    mem[16'h149C] = 8'h00;
    mem[16'h149D] = 8'h00;
    mem[16'h149E] = 8'h04; // PUSH RAX
    mem[16'h149F] = 8'h00;
    mem[16'h14A0] = 8'h85; // SUBN RSP 8
    mem[16'h14A1] = 8'h06;
    mem[16'h14A2] = 8'h08;
    mem[16'h14A3] = 8'h00;
    mem[16'h14A4] = 8'h00;
    mem[16'h14A5] = 8'h00;
    mem[16'h14A6] = 8'h05; // PUSHN 1
    mem[16'h14A7] = 8'h00;
    mem[16'h14A8] = 8'h01;
    mem[16'h14A9] = 8'h00;
    mem[16'h14AA] = 8'h00;
    mem[16'h14AB] = 8'h00;
    mem[16'h14AC] = 8'h08; // POP RDI
    mem[16'h14AD] = 8'h01;
    mem[16'h14AE] = 8'h81; // ADDN RSP 8
    mem[16'h14AF] = 8'h06;
    mem[16'h14B0] = 8'h08;
    mem[16'h14B1] = 8'h00;
    mem[16'h14B2] = 8'h00;
    mem[16'h14B3] = 8'h00;
    mem[16'h14B4] = 8'h08; // POP RAX
    mem[16'h14B5] = 8'h00;
    mem[16'h14B6] = 8'h81; // ADDN RSP 8
    mem[16'h14B7] = 8'h06;
    mem[16'h14B8] = 8'h08;
    mem[16'h14B9] = 8'h00;
    mem[16'h14BA] = 8'h00;
    mem[16'h14BB] = 8'h00;
    mem[16'h14BC] = 8'h80; // ADD RAX RDI
    mem[16'h14BD] = 8'h00;
    mem[16'h14BE] = 8'h01;
    mem[16'h14BF] = 8'h85; // SUBN RSP 8
    mem[16'h14C0] = 8'h06;
    mem[16'h14C1] = 8'h08;
    mem[16'h14C2] = 8'h00;
    mem[16'h14C3] = 8'h00;
    mem[16'h14C4] = 8'h00;
    mem[16'h14C5] = 8'h04; // PUSH RAX
    mem[16'h14C6] = 8'h00;
    mem[16'h14C7] = 8'h08; // POP RDI
    mem[16'h14C8] = 8'h01;
    mem[16'h14C9] = 8'h81; // ADDN RSP 8
    mem[16'h14CA] = 8'h06;
    mem[16'h14CB] = 8'h08;
    mem[16'h14CC] = 8'h00;
    mem[16'h14CD] = 8'h00;
    mem[16'h14CE] = 8'h00;
    mem[16'h14CF] = 8'h08; // POP RAX
    mem[16'h14D0] = 8'h00;
    mem[16'h14D1] = 8'h81; // ADDN RSP 8
    mem[16'h14D2] = 8'h06;
    mem[16'h14D3] = 8'h08;
    mem[16'h14D4] = 8'h00;
    mem[16'h14D5] = 8'h00;
    mem[16'h14D6] = 8'h00;
    mem[16'h14D7] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h14D8] = 8'h00;
    mem[16'h14D9] = 8'h01;
    mem[16'h14DA] = 8'h85; // SUBN RSP 8
    mem[16'h14DB] = 8'h06;
    mem[16'h14DC] = 8'h08;
    mem[16'h14DD] = 8'h00;
    mem[16'h14DE] = 8'h00;
    mem[16'h14DF] = 8'h00;
    mem[16'h14E0] = 8'h04; // PUSH RDI
    mem[16'h14E1] = 8'h01;
    mem[16'h14E2] = 8'h81; // ADDN RSP 8
    mem[16'h14E3] = 8'h06;
    mem[16'h14E4] = 8'h08;
    mem[16'h14E5] = 8'h00;
    mem[16'h14E6] = 8'h00;
    mem[16'h14E7] = 8'h00;
    mem[16'h14E8] = 8'h40; // MOV RAX RBP
    mem[16'h14E9] = 8'h00;
    mem[16'h14EA] = 8'h05;
    mem[16'h14EB] = 8'h85; // SUBN RAX 12
    mem[16'h14EC] = 8'h00;
    mem[16'h14ED] = 8'h0C;
    mem[16'h14EE] = 8'h00;
    mem[16'h14EF] = 8'h00;
    mem[16'h14F0] = 8'h00;
    mem[16'h14F1] = 8'h85; // SUBN RSP 8
    mem[16'h14F2] = 8'h06;
    mem[16'h14F3] = 8'h08;
    mem[16'h14F4] = 8'h00;
    mem[16'h14F5] = 8'h00;
    mem[16'h14F6] = 8'h00;
    mem[16'h14F7] = 8'h04; // PUSH RAX
    mem[16'h14F8] = 8'h00;
    mem[16'h14F9] = 8'h40; // MOV RAX RBP
    mem[16'h14FA] = 8'h00;
    mem[16'h14FB] = 8'h05;
    mem[16'h14FC] = 8'h85; // SUBN RAX 12
    mem[16'h14FD] = 8'h00;
    mem[16'h14FE] = 8'h0C;
    mem[16'h14FF] = 8'h00;
    mem[16'h1500] = 8'h00;
    mem[16'h1501] = 8'h00;
    mem[16'h1502] = 8'h85; // SUBN RSP 8
    mem[16'h1503] = 8'h06;
    mem[16'h1504] = 8'h08;
    mem[16'h1505] = 8'h00;
    mem[16'h1506] = 8'h00;
    mem[16'h1507] = 8'h00;
    mem[16'h1508] = 8'h04; // PUSH RAX
    mem[16'h1509] = 8'h00;
    mem[16'h150A] = 8'h08; // POP RAX
    mem[16'h150B] = 8'h00;
    mem[16'h150C] = 8'h81; // ADDN RSP 8
    mem[16'h150D] = 8'h06;
    mem[16'h150E] = 8'h08;
    mem[16'h150F] = 8'h00;
    mem[16'h1510] = 8'h00;
    mem[16'h1511] = 8'h00;
    mem[16'h1512] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1513] = 8'h00;
    mem[16'h1514] = 8'h00;
    mem[16'h1515] = 8'h85; // SUBN RSP 8
    mem[16'h1516] = 8'h06;
    mem[16'h1517] = 8'h08;
    mem[16'h1518] = 8'h00;
    mem[16'h1519] = 8'h00;
    mem[16'h151A] = 8'h00;
    mem[16'h151B] = 8'h04; // PUSH RAX
    mem[16'h151C] = 8'h00;
    mem[16'h151D] = 8'h85; // SUBN RSP 8
    mem[16'h151E] = 8'h06;
    mem[16'h151F] = 8'h08;
    mem[16'h1520] = 8'h00;
    mem[16'h1521] = 8'h00;
    mem[16'h1522] = 8'h00;
    mem[16'h1523] = 8'h05; // PUSHN 1
    mem[16'h1524] = 8'h00;
    mem[16'h1525] = 8'h01;
    mem[16'h1526] = 8'h00;
    mem[16'h1527] = 8'h00;
    mem[16'h1528] = 8'h00;
    mem[16'h1529] = 8'h08; // POP RDI
    mem[16'h152A] = 8'h01;
    mem[16'h152B] = 8'h81; // ADDN RSP 8
    mem[16'h152C] = 8'h06;
    mem[16'h152D] = 8'h08;
    mem[16'h152E] = 8'h00;
    mem[16'h152F] = 8'h00;
    mem[16'h1530] = 8'h00;
    mem[16'h1531] = 8'h08; // POP RAX
    mem[16'h1532] = 8'h00;
    mem[16'h1533] = 8'h81; // ADDN RSP 8
    mem[16'h1534] = 8'h06;
    mem[16'h1535] = 8'h08;
    mem[16'h1536] = 8'h00;
    mem[16'h1537] = 8'h00;
    mem[16'h1538] = 8'h00;
    mem[16'h1539] = 8'h84; // SUB RAX RDI
    mem[16'h153A] = 8'h00;
    mem[16'h153B] = 8'h01;
    mem[16'h153C] = 8'h85; // SUBN RSP 8
    mem[16'h153D] = 8'h06;
    mem[16'h153E] = 8'h08;
    mem[16'h153F] = 8'h00;
    mem[16'h1540] = 8'h00;
    mem[16'h1541] = 8'h00;
    mem[16'h1542] = 8'h04; // PUSH RAX
    mem[16'h1543] = 8'h00;
    mem[16'h1544] = 8'h08; // POP RDI
    mem[16'h1545] = 8'h01;
    mem[16'h1546] = 8'h81; // ADDN RSP 8
    mem[16'h1547] = 8'h06;
    mem[16'h1548] = 8'h08;
    mem[16'h1549] = 8'h00;
    mem[16'h154A] = 8'h00;
    mem[16'h154B] = 8'h00;
    mem[16'h154C] = 8'h08; // POP RAX
    mem[16'h154D] = 8'h00;
    mem[16'h154E] = 8'h81; // ADDN RSP 8
    mem[16'h154F] = 8'h06;
    mem[16'h1550] = 8'h08;
    mem[16'h1551] = 8'h00;
    mem[16'h1552] = 8'h00;
    mem[16'h1553] = 8'h00;
    mem[16'h1554] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h1555] = 8'h00;
    mem[16'h1556] = 8'h01;
    mem[16'h1557] = 8'h85; // SUBN RSP 8
    mem[16'h1558] = 8'h06;
    mem[16'h1559] = 8'h08;
    mem[16'h155A] = 8'h00;
    mem[16'h155B] = 8'h00;
    mem[16'h155C] = 8'h00;
    mem[16'h155D] = 8'h04; // PUSH RDI
    mem[16'h155E] = 8'h01;
    mem[16'h155F] = 8'h81; // ADDN RSP 8
    mem[16'h1560] = 8'h06;
    mem[16'h1561] = 8'h08;
    mem[16'h1562] = 8'h00;
    mem[16'h1563] = 8'h00;
    mem[16'h1564] = 8'h00;
    mem[16'h1565] = 8'h40; // MOV RAX RBP
    mem[16'h1566] = 8'h00;
    mem[16'h1567] = 8'h05;
    mem[16'h1568] = 8'h85; // SUBN RAX 4
    mem[16'h1569] = 8'h00;
    mem[16'h156A] = 8'h04;
    mem[16'h156B] = 8'h00;
    mem[16'h156C] = 8'h00;
    mem[16'h156D] = 8'h00;
    mem[16'h156E] = 8'h85; // SUBN RSP 8
    mem[16'h156F] = 8'h06;
    mem[16'h1570] = 8'h08;
    mem[16'h1571] = 8'h00;
    mem[16'h1572] = 8'h00;
    mem[16'h1573] = 8'h00;
    mem[16'h1574] = 8'h04; // PUSH RAX
    mem[16'h1575] = 8'h00;
    mem[16'h1576] = 8'h40; // MOV RAX RBP
    mem[16'h1577] = 8'h00;
    mem[16'h1578] = 8'h05;
    mem[16'h1579] = 8'h85; // SUBN RAX 4
    mem[16'h157A] = 8'h00;
    mem[16'h157B] = 8'h04;
    mem[16'h157C] = 8'h00;
    mem[16'h157D] = 8'h00;
    mem[16'h157E] = 8'h00;
    mem[16'h157F] = 8'h85; // SUBN RSP 8
    mem[16'h1580] = 8'h06;
    mem[16'h1581] = 8'h08;
    mem[16'h1582] = 8'h00;
    mem[16'h1583] = 8'h00;
    mem[16'h1584] = 8'h00;
    mem[16'h1585] = 8'h04; // PUSH RAX
    mem[16'h1586] = 8'h00;
    mem[16'h1587] = 8'h08; // POP RAX
    mem[16'h1588] = 8'h00;
    mem[16'h1589] = 8'h81; // ADDN RSP 8
    mem[16'h158A] = 8'h06;
    mem[16'h158B] = 8'h08;
    mem[16'h158C] = 8'h00;
    mem[16'h158D] = 8'h00;
    mem[16'h158E] = 8'h00;
    mem[16'h158F] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1590] = 8'h00;
    mem[16'h1591] = 8'h00;
    mem[16'h1592] = 8'h85; // SUBN RSP 8
    mem[16'h1593] = 8'h06;
    mem[16'h1594] = 8'h08;
    mem[16'h1595] = 8'h00;
    mem[16'h1596] = 8'h00;
    mem[16'h1597] = 8'h00;
    mem[16'h1598] = 8'h04; // PUSH RAX
    mem[16'h1599] = 8'h00;
    mem[16'h159A] = 8'h85; // SUBN RSP 8
    mem[16'h159B] = 8'h06;
    mem[16'h159C] = 8'h08;
    mem[16'h159D] = 8'h00;
    mem[16'h159E] = 8'h00;
    mem[16'h159F] = 8'h00;
    mem[16'h15A0] = 8'h05; // PUSHN 1
    mem[16'h15A1] = 8'h00;
    mem[16'h15A2] = 8'h01;
    mem[16'h15A3] = 8'h00;
    mem[16'h15A4] = 8'h00;
    mem[16'h15A5] = 8'h00;
    mem[16'h15A6] = 8'h08; // POP RDI
    mem[16'h15A7] = 8'h01;
    mem[16'h15A8] = 8'h81; // ADDN RSP 8
    mem[16'h15A9] = 8'h06;
    mem[16'h15AA] = 8'h08;
    mem[16'h15AB] = 8'h00;
    mem[16'h15AC] = 8'h00;
    mem[16'h15AD] = 8'h00;
    mem[16'h15AE] = 8'h08; // POP RAX
    mem[16'h15AF] = 8'h00;
    mem[16'h15B0] = 8'h81; // ADDN RSP 8
    mem[16'h15B1] = 8'h06;
    mem[16'h15B2] = 8'h08;
    mem[16'h15B3] = 8'h00;
    mem[16'h15B4] = 8'h00;
    mem[16'h15B5] = 8'h00;
    mem[16'h15B6] = 8'h80; // ADD RAX RDI
    mem[16'h15B7] = 8'h00;
    mem[16'h15B8] = 8'h01;
    mem[16'h15B9] = 8'h85; // SUBN RSP 8
    mem[16'h15BA] = 8'h06;
    mem[16'h15BB] = 8'h08;
    mem[16'h15BC] = 8'h00;
    mem[16'h15BD] = 8'h00;
    mem[16'h15BE] = 8'h00;
    mem[16'h15BF] = 8'h04; // PUSH RAX
    mem[16'h15C0] = 8'h00;
    mem[16'h15C1] = 8'h08; // POP RDI
    mem[16'h15C2] = 8'h01;
    mem[16'h15C3] = 8'h81; // ADDN RSP 8
    mem[16'h15C4] = 8'h06;
    mem[16'h15C5] = 8'h08;
    mem[16'h15C6] = 8'h00;
    mem[16'h15C7] = 8'h00;
    mem[16'h15C8] = 8'h00;
    mem[16'h15C9] = 8'h08; // POP RAX
    mem[16'h15CA] = 8'h00;
    mem[16'h15CB] = 8'h81; // ADDN RSP 8
    mem[16'h15CC] = 8'h06;
    mem[16'h15CD] = 8'h08;
    mem[16'h15CE] = 8'h00;
    mem[16'h15CF] = 8'h00;
    mem[16'h15D0] = 8'h00;
    mem[16'h15D1] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h15D2] = 8'h00;
    mem[16'h15D3] = 8'h01;
    mem[16'h15D4] = 8'h85; // SUBN RSP 8
    mem[16'h15D5] = 8'h06;
    mem[16'h15D6] = 8'h08;
    mem[16'h15D7] = 8'h00;
    mem[16'h15D8] = 8'h00;
    mem[16'h15D9] = 8'h00;
    mem[16'h15DA] = 8'h04; // PUSH RDI
    mem[16'h15DB] = 8'h01;
    mem[16'h15DC] = 8'h81; // ADDN RSP 8
    mem[16'h15DD] = 8'h06;
    mem[16'h15DE] = 8'h08;
    mem[16'h15DF] = 8'h00;
    mem[16'h15E0] = 8'h00;
    mem[16'h15E1] = 8'h00;
    mem[16'h15E2] = 8'h22; // JMP .Lbegin9
    mem[16'h15E3] = 8'hAE;
    mem[16'h15E4] = 8'h10;
    mem[16'h15E5] = 8'h00;
    mem[16'h15E6] = 8'h00;
    mem[16'h15E7] = 8'h00;
    mem[16'h15E8] = 8'h00;
    mem[16'h15E9] = 8'h00;
    mem[16'h15EA] = 8'h00;
                          // .Lend9:
    mem[16'h15EB] = 8'h85; // SUBN RSP 8
    mem[16'h15EC] = 8'h06;
    mem[16'h15ED] = 8'h08;
    mem[16'h15EE] = 8'h00;
    mem[16'h15EF] = 8'h00;
    mem[16'h15F0] = 8'h00;
    mem[16'h15F1] = 8'h05; // PUSHN 1
    mem[16'h15F2] = 8'h00;
    mem[16'h15F3] = 8'h01;
    mem[16'h15F4] = 8'h00;
    mem[16'h15F5] = 8'h00;
    mem[16'h15F6] = 8'h00;
    mem[16'h15F7] = 8'h08; // POP RAX
    mem[16'h15F8] = 8'h00;
    mem[16'h15F9] = 8'h81; // ADDN RSP 8
    mem[16'h15FA] = 8'h06;
    mem[16'h15FB] = 8'h08;
    mem[16'h15FC] = 8'h00;
    mem[16'h15FD] = 8'h00;
    mem[16'h15FE] = 8'h00;
    mem[16'h15FF] = 8'h22; // JMP .Lreturn.check
    mem[16'h1600] = 8'h08;
    mem[16'h1601] = 8'h16;
    mem[16'h1602] = 8'h00;
    mem[16'h1603] = 8'h00;
    mem[16'h1604] = 8'h00;
    mem[16'h1605] = 8'h00;
    mem[16'h1606] = 8'h00;
    mem[16'h1607] = 8'h00;
                          // .Lreturn.check:
    mem[16'h1608] = 8'h40; // MOV RSP RBP
    mem[16'h1609] = 8'h06;
    mem[16'h160A] = 8'h05;
    mem[16'h160B] = 8'h08; // POP RBP
    mem[16'h160C] = 8'h05;
    mem[16'h160D] = 8'h81; // ADDN RSP 8
    mem[16'h160E] = 8'h06;
    mem[16'h160F] = 8'h08;
    mem[16'h1610] = 8'h00;
    mem[16'h1611] = 8'h00;
    mem[16'h1612] = 8'h00;
    mem[16'h1613] = 8'h08; // POP RBX
    mem[16'h1614] = 8'h07;
    mem[16'h1615] = 8'h81; // ADDN RSP 8
    mem[16'h1616] = 8'h06;
    mem[16'h1617] = 8'h08;
    mem[16'h1618] = 8'h00;
    mem[16'h1619] = 8'h00;
    mem[16'h161A] = 8'h00;
    mem[16'h161B] = 8'h20; // JMPR RBX
    mem[16'h161C] = 8'h07;
                          // eightqueen:
    mem[16'h161D] = 8'h85; // SUBN RSP 8
    mem[16'h161E] = 8'h06;
    mem[16'h161F] = 8'h08;
    mem[16'h1620] = 8'h00;
    mem[16'h1621] = 8'h00;
    mem[16'h1622] = 8'h00;
    mem[16'h1623] = 8'h04; // PUSH RBP
    mem[16'h1624] = 8'h05;
    mem[16'h1625] = 8'h40; // MOV RBP RSP
    mem[16'h1626] = 8'h05;
    mem[16'h1627] = 8'h06;
    mem[16'h1628] = 8'h85; // SUBN RSP 16
    mem[16'h1629] = 8'h06;
    mem[16'h162A] = 8'h10;
    mem[16'h162B] = 8'h00;
    mem[16'h162C] = 8'h00;
    mem[16'h162D] = 8'h00;
    mem[16'h162E] = 8'h40; // MOV RBX RBP
    mem[16'h162F] = 8'h07;
    mem[16'h1630] = 8'h05;
    mem[16'h1631] = 8'h85; // SUBN RBX 12
    mem[16'h1632] = 8'h07;
    mem[16'h1633] = 8'h0C;
    mem[16'h1634] = 8'h00;
    mem[16'h1635] = 8'h00;
    mem[16'h1636] = 8'h00;
    mem[16'h1637] = 8'h58; // MOVAR4 RBX RDI
    mem[16'h1638] = 8'h07;
    mem[16'h1639] = 8'h01;
    mem[16'h163A] = 8'h40; // MOV RAX RBP
    mem[16'h163B] = 8'h00;
    mem[16'h163C] = 8'h05;
    mem[16'h163D] = 8'h85; // SUBN RAX 12
    mem[16'h163E] = 8'h00;
    mem[16'h163F] = 8'h0C;
    mem[16'h1640] = 8'h00;
    mem[16'h1641] = 8'h00;
    mem[16'h1642] = 8'h00;
    mem[16'h1643] = 8'h85; // SUBN RSP 8
    mem[16'h1644] = 8'h06;
    mem[16'h1645] = 8'h08;
    mem[16'h1646] = 8'h00;
    mem[16'h1647] = 8'h00;
    mem[16'h1648] = 8'h00;
    mem[16'h1649] = 8'h04; // PUSH RAX
    mem[16'h164A] = 8'h00;
    mem[16'h164B] = 8'h08; // POP RAX
    mem[16'h164C] = 8'h00;
    mem[16'h164D] = 8'h81; // ADDN RSP 8
    mem[16'h164E] = 8'h06;
    mem[16'h164F] = 8'h08;
    mem[16'h1650] = 8'h00;
    mem[16'h1651] = 8'h00;
    mem[16'h1652] = 8'h00;
    mem[16'h1653] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1654] = 8'h00;
    mem[16'h1655] = 8'h00;
    mem[16'h1656] = 8'h85; // SUBN RSP 8
    mem[16'h1657] = 8'h06;
    mem[16'h1658] = 8'h08;
    mem[16'h1659] = 8'h00;
    mem[16'h165A] = 8'h00;
    mem[16'h165B] = 8'h00;
    mem[16'h165C] = 8'h04; // PUSH RAX
    mem[16'h165D] = 8'h00;
    mem[16'h165E] = 8'h85; // SUBN RSP 8
    mem[16'h165F] = 8'h06;
    mem[16'h1660] = 8'h08;
    mem[16'h1661] = 8'h00;
    mem[16'h1662] = 8'h00;
    mem[16'h1663] = 8'h00;
    mem[16'h1664] = 8'h05; // PUSHN 8
    mem[16'h1665] = 8'h00;
    mem[16'h1666] = 8'h08;
    mem[16'h1667] = 8'h00;
    mem[16'h1668] = 8'h00;
    mem[16'h1669] = 8'h00;
    mem[16'h166A] = 8'h08; // POP RDI
    mem[16'h166B] = 8'h01;
    mem[16'h166C] = 8'h81; // ADDN RSP 8
    mem[16'h166D] = 8'h06;
    mem[16'h166E] = 8'h08;
    mem[16'h166F] = 8'h00;
    mem[16'h1670] = 8'h00;
    mem[16'h1671] = 8'h00;
    mem[16'h1672] = 8'h08; // POP RAX
    mem[16'h1673] = 8'h00;
    mem[16'h1674] = 8'h81; // ADDN RSP 8
    mem[16'h1675] = 8'h06;
    mem[16'h1676] = 8'h08;
    mem[16'h1677] = 8'h00;
    mem[16'h1678] = 8'h00;
    mem[16'h1679] = 8'h00;
    mem[16'h167A] = 8'h90; // CMP RAX RDI
    mem[16'h167B] = 8'h00;
    mem[16'h167C] = 8'h01;
    mem[16'h167D] = 8'h10; // SETE RAX
    mem[16'h167E] = 8'h00;
    mem[16'h167F] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h1680] = 8'h00;
    mem[16'h1681] = 8'h00;
    mem[16'h1682] = 8'h85; // SUBN RSP 8
    mem[16'h1683] = 8'h06;
    mem[16'h1684] = 8'h08;
    mem[16'h1685] = 8'h00;
    mem[16'h1686] = 8'h00;
    mem[16'h1687] = 8'h00;
    mem[16'h1688] = 8'h04; // PUSH RAX
    mem[16'h1689] = 8'h00;
    mem[16'h168A] = 8'h08; // POP RAX
    mem[16'h168B] = 8'h00;
    mem[16'h168C] = 8'h81; // ADDN RSP 8
    mem[16'h168D] = 8'h06;
    mem[16'h168E] = 8'h08;
    mem[16'h168F] = 8'h00;
    mem[16'h1690] = 8'h00;
    mem[16'h1691] = 8'h00;
    mem[16'h1692] = 8'h91; // CMPN RAX 0
    mem[16'h1693] = 8'h00;
    mem[16'h1694] = 8'h00;
    mem[16'h1695] = 8'h00;
    mem[16'h1696] = 8'h00;
    mem[16'h1697] = 8'h00;
    mem[16'h1698] = 8'h26; // JE .Lend13
    mem[16'h1699] = 8'hBE;
    mem[16'h169A] = 8'h16;
    mem[16'h169B] = 8'h00;
    mem[16'h169C] = 8'h00;
    mem[16'h169D] = 8'h00;
    mem[16'h169E] = 8'h00;
    mem[16'h169F] = 8'h00;
    mem[16'h16A0] = 8'h00;
    mem[16'h16A1] = 8'h85; // SUBN RSP 8
    mem[16'h16A2] = 8'h06;
    mem[16'h16A3] = 8'h08;
    mem[16'h16A4] = 8'h00;
    mem[16'h16A5] = 8'h00;
    mem[16'h16A6] = 8'h00;
    mem[16'h16A7] = 8'h05; // PUSHN 1
    mem[16'h16A8] = 8'h00;
    mem[16'h16A9] = 8'h01;
    mem[16'h16AA] = 8'h00;
    mem[16'h16AB] = 8'h00;
    mem[16'h16AC] = 8'h00;
    mem[16'h16AD] = 8'h08; // POP RAX
    mem[16'h16AE] = 8'h00;
    mem[16'h16AF] = 8'h81; // ADDN RSP 8
    mem[16'h16B0] = 8'h06;
    mem[16'h16B1] = 8'h08;
    mem[16'h16B2] = 8'h00;
    mem[16'h16B3] = 8'h00;
    mem[16'h16B4] = 8'h00;
    mem[16'h16B5] = 8'h22; // JMP .Lreturn.eightqueen
    mem[16'h16B6] = 8'hB9;
    mem[16'h16B7] = 8'h1C;
    mem[16'h16B8] = 8'h00;
    mem[16'h16B9] = 8'h00;
    mem[16'h16BA] = 8'h00;
    mem[16'h16BB] = 8'h00;
    mem[16'h16BC] = 8'h00;
    mem[16'h16BD] = 8'h00;
                          // .Lend13:
    mem[16'h16BE] = 8'h40; // MOV RAX RBP
    mem[16'h16BF] = 8'h00;
    mem[16'h16C0] = 8'h05;
    mem[16'h16C1] = 8'h85; // SUBN RAX 4
    mem[16'h16C2] = 8'h00;
    mem[16'h16C3] = 8'h04;
    mem[16'h16C4] = 8'h00;
    mem[16'h16C5] = 8'h00;
    mem[16'h16C6] = 8'h00;
    mem[16'h16C7] = 8'h85; // SUBN RSP 8
    mem[16'h16C8] = 8'h06;
    mem[16'h16C9] = 8'h08;
    mem[16'h16CA] = 8'h00;
    mem[16'h16CB] = 8'h00;
    mem[16'h16CC] = 8'h00;
    mem[16'h16CD] = 8'h04; // PUSH RAX
    mem[16'h16CE] = 8'h00;
    mem[16'h16CF] = 8'h85; // SUBN RSP 8
    mem[16'h16D0] = 8'h06;
    mem[16'h16D1] = 8'h08;
    mem[16'h16D2] = 8'h00;
    mem[16'h16D3] = 8'h00;
    mem[16'h16D4] = 8'h00;
    mem[16'h16D5] = 8'h05; // PUSHN 0
    mem[16'h16D6] = 8'h00;
    mem[16'h16D7] = 8'h00;
    mem[16'h16D8] = 8'h00;
    mem[16'h16D9] = 8'h00;
    mem[16'h16DA] = 8'h00;
    mem[16'h16DB] = 8'h08; // POP RDI
    mem[16'h16DC] = 8'h01;
    mem[16'h16DD] = 8'h81; // ADDN RSP 8
    mem[16'h16DE] = 8'h06;
    mem[16'h16DF] = 8'h08;
    mem[16'h16E0] = 8'h00;
    mem[16'h16E1] = 8'h00;
    mem[16'h16E2] = 8'h00;
    mem[16'h16E3] = 8'h08; // POP RAX
    mem[16'h16E4] = 8'h00;
    mem[16'h16E5] = 8'h81; // ADDN RSP 8
    mem[16'h16E6] = 8'h06;
    mem[16'h16E7] = 8'h08;
    mem[16'h16E8] = 8'h00;
    mem[16'h16E9] = 8'h00;
    mem[16'h16EA] = 8'h00;
    mem[16'h16EB] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h16EC] = 8'h00;
    mem[16'h16ED] = 8'h01;
    mem[16'h16EE] = 8'h85; // SUBN RSP 8
    mem[16'h16EF] = 8'h06;
    mem[16'h16F0] = 8'h08;
    mem[16'h16F1] = 8'h00;
    mem[16'h16F2] = 8'h00;
    mem[16'h16F3] = 8'h00;
    mem[16'h16F4] = 8'h04; // PUSH RDI
    mem[16'h16F5] = 8'h01;
    mem[16'h16F6] = 8'h81; // ADDN RSP 8
    mem[16'h16F7] = 8'h06;
    mem[16'h16F8] = 8'h08;
    mem[16'h16F9] = 8'h00;
    mem[16'h16FA] = 8'h00;
    mem[16'h16FB] = 8'h00;
                          // .Lbegin14:
    mem[16'h16FC] = 8'h40; // MOV RAX RBP
    mem[16'h16FD] = 8'h00;
    mem[16'h16FE] = 8'h05;
    mem[16'h16FF] = 8'h85; // SUBN RAX 4
    mem[16'h1700] = 8'h00;
    mem[16'h1701] = 8'h04;
    mem[16'h1702] = 8'h00;
    mem[16'h1703] = 8'h00;
    mem[16'h1704] = 8'h00;
    mem[16'h1705] = 8'h85; // SUBN RSP 8
    mem[16'h1706] = 8'h06;
    mem[16'h1707] = 8'h08;
    mem[16'h1708] = 8'h00;
    mem[16'h1709] = 8'h00;
    mem[16'h170A] = 8'h00;
    mem[16'h170B] = 8'h04; // PUSH RAX
    mem[16'h170C] = 8'h00;
    mem[16'h170D] = 8'h08; // POP RAX
    mem[16'h170E] = 8'h00;
    mem[16'h170F] = 8'h81; // ADDN RSP 8
    mem[16'h1710] = 8'h06;
    mem[16'h1711] = 8'h08;
    mem[16'h1712] = 8'h00;
    mem[16'h1713] = 8'h00;
    mem[16'h1714] = 8'h00;
    mem[16'h1715] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1716] = 8'h00;
    mem[16'h1717] = 8'h00;
    mem[16'h1718] = 8'h85; // SUBN RSP 8
    mem[16'h1719] = 8'h06;
    mem[16'h171A] = 8'h08;
    mem[16'h171B] = 8'h00;
    mem[16'h171C] = 8'h00;
    mem[16'h171D] = 8'h00;
    mem[16'h171E] = 8'h04; // PUSH RAX
    mem[16'h171F] = 8'h00;
    mem[16'h1720] = 8'h85; // SUBN RSP 8
    mem[16'h1721] = 8'h06;
    mem[16'h1722] = 8'h08;
    mem[16'h1723] = 8'h00;
    mem[16'h1724] = 8'h00;
    mem[16'h1725] = 8'h00;
    mem[16'h1726] = 8'h05; // PUSHN 8
    mem[16'h1727] = 8'h00;
    mem[16'h1728] = 8'h08;
    mem[16'h1729] = 8'h00;
    mem[16'h172A] = 8'h00;
    mem[16'h172B] = 8'h00;
    mem[16'h172C] = 8'h08; // POP RDI
    mem[16'h172D] = 8'h01;
    mem[16'h172E] = 8'h81; // ADDN RSP 8
    mem[16'h172F] = 8'h06;
    mem[16'h1730] = 8'h08;
    mem[16'h1731] = 8'h00;
    mem[16'h1732] = 8'h00;
    mem[16'h1733] = 8'h00;
    mem[16'h1734] = 8'h08; // POP RAX
    mem[16'h1735] = 8'h00;
    mem[16'h1736] = 8'h81; // ADDN RSP 8
    mem[16'h1737] = 8'h06;
    mem[16'h1738] = 8'h08;
    mem[16'h1739] = 8'h00;
    mem[16'h173A] = 8'h00;
    mem[16'h173B] = 8'h00;
    mem[16'h173C] = 8'h90; // CMP RAX RDI
    mem[16'h173D] = 8'h00;
    mem[16'h173E] = 8'h01;
    mem[16'h173F] = 8'h18; // SETL RAX
    mem[16'h1740] = 8'h00;
    mem[16'h1741] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h1742] = 8'h00;
    mem[16'h1743] = 8'h00;
    mem[16'h1744] = 8'h85; // SUBN RSP 8
    mem[16'h1745] = 8'h06;
    mem[16'h1746] = 8'h08;
    mem[16'h1747] = 8'h00;
    mem[16'h1748] = 8'h00;
    mem[16'h1749] = 8'h00;
    mem[16'h174A] = 8'h04; // PUSH RAX
    mem[16'h174B] = 8'h00;
    mem[16'h174C] = 8'h08; // POP RAX
    mem[16'h174D] = 8'h00;
    mem[16'h174E] = 8'h81; // ADDN RSP 8
    mem[16'h174F] = 8'h06;
    mem[16'h1750] = 8'h08;
    mem[16'h1751] = 8'h00;
    mem[16'h1752] = 8'h00;
    mem[16'h1753] = 8'h00;
    mem[16'h1754] = 8'h91; // CMPN RAX 0
    mem[16'h1755] = 8'h00;
    mem[16'h1756] = 8'h00;
    mem[16'h1757] = 8'h00;
    mem[16'h1758] = 8'h00;
    mem[16'h1759] = 8'h00;
    mem[16'h175A] = 8'h26; // JE .Lend14
    mem[16'h175B] = 8'h9C;
    mem[16'h175C] = 8'h1C;
    mem[16'h175D] = 8'h00;
    mem[16'h175E] = 8'h00;
    mem[16'h175F] = 8'h00;
    mem[16'h1760] = 8'h00;
    mem[16'h1761] = 8'h00;
    mem[16'h1762] = 8'h00;
    mem[16'h1763] = 8'h40; // MOV RAX RBP
    mem[16'h1764] = 8'h00;
    mem[16'h1765] = 8'h05;
    mem[16'h1766] = 8'h85; // SUBN RAX 8
    mem[16'h1767] = 8'h00;
    mem[16'h1768] = 8'h08;
    mem[16'h1769] = 8'h00;
    mem[16'h176A] = 8'h00;
    mem[16'h176B] = 8'h00;
    mem[16'h176C] = 8'h85; // SUBN RSP 8
    mem[16'h176D] = 8'h06;
    mem[16'h176E] = 8'h08;
    mem[16'h176F] = 8'h00;
    mem[16'h1770] = 8'h00;
    mem[16'h1771] = 8'h00;
    mem[16'h1772] = 8'h04; // PUSH RAX
    mem[16'h1773] = 8'h00;
    mem[16'h1774] = 8'h85; // SUBN RSP 8
    mem[16'h1775] = 8'h06;
    mem[16'h1776] = 8'h08;
    mem[16'h1777] = 8'h00;
    mem[16'h1778] = 8'h00;
    mem[16'h1779] = 8'h00;
    mem[16'h177A] = 8'h05; // PUSHN 0
    mem[16'h177B] = 8'h00;
    mem[16'h177C] = 8'h00;
    mem[16'h177D] = 8'h00;
    mem[16'h177E] = 8'h00;
    mem[16'h177F] = 8'h00;
    mem[16'h1780] = 8'h08; // POP RDI
    mem[16'h1781] = 8'h01;
    mem[16'h1782] = 8'h81; // ADDN RSP 8
    mem[16'h1783] = 8'h06;
    mem[16'h1784] = 8'h08;
    mem[16'h1785] = 8'h00;
    mem[16'h1786] = 8'h00;
    mem[16'h1787] = 8'h00;
    mem[16'h1788] = 8'h08; // POP RAX
    mem[16'h1789] = 8'h00;
    mem[16'h178A] = 8'h81; // ADDN RSP 8
    mem[16'h178B] = 8'h06;
    mem[16'h178C] = 8'h08;
    mem[16'h178D] = 8'h00;
    mem[16'h178E] = 8'h00;
    mem[16'h178F] = 8'h00;
    mem[16'h1790] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h1791] = 8'h00;
    mem[16'h1792] = 8'h01;
    mem[16'h1793] = 8'h85; // SUBN RSP 8
    mem[16'h1794] = 8'h06;
    mem[16'h1795] = 8'h08;
    mem[16'h1796] = 8'h00;
    mem[16'h1797] = 8'h00;
    mem[16'h1798] = 8'h00;
    mem[16'h1799] = 8'h04; // PUSH RDI
    mem[16'h179A] = 8'h01;
    mem[16'h179B] = 8'h81; // ADDN RSP 8
    mem[16'h179C] = 8'h06;
    mem[16'h179D] = 8'h08;
    mem[16'h179E] = 8'h00;
    mem[16'h179F] = 8'h00;
    mem[16'h17A0] = 8'h00;
                          // .Lbegin15:
    mem[16'h17A1] = 8'h40; // MOV RAX RBP
    mem[16'h17A2] = 8'h00;
    mem[16'h17A3] = 8'h05;
    mem[16'h17A4] = 8'h85; // SUBN RAX 8
    mem[16'h17A5] = 8'h00;
    mem[16'h17A6] = 8'h08;
    mem[16'h17A7] = 8'h00;
    mem[16'h17A8] = 8'h00;
    mem[16'h17A9] = 8'h00;
    mem[16'h17AA] = 8'h85; // SUBN RSP 8
    mem[16'h17AB] = 8'h06;
    mem[16'h17AC] = 8'h08;
    mem[16'h17AD] = 8'h00;
    mem[16'h17AE] = 8'h00;
    mem[16'h17AF] = 8'h00;
    mem[16'h17B0] = 8'h04; // PUSH RAX
    mem[16'h17B1] = 8'h00;
    mem[16'h17B2] = 8'h08; // POP RAX
    mem[16'h17B3] = 8'h00;
    mem[16'h17B4] = 8'h81; // ADDN RSP 8
    mem[16'h17B5] = 8'h06;
    mem[16'h17B6] = 8'h08;
    mem[16'h17B7] = 8'h00;
    mem[16'h17B8] = 8'h00;
    mem[16'h17B9] = 8'h00;
    mem[16'h17BA] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h17BB] = 8'h00;
    mem[16'h17BC] = 8'h00;
    mem[16'h17BD] = 8'h85; // SUBN RSP 8
    mem[16'h17BE] = 8'h06;
    mem[16'h17BF] = 8'h08;
    mem[16'h17C0] = 8'h00;
    mem[16'h17C1] = 8'h00;
    mem[16'h17C2] = 8'h00;
    mem[16'h17C3] = 8'h04; // PUSH RAX
    mem[16'h17C4] = 8'h00;
    mem[16'h17C5] = 8'h85; // SUBN RSP 8
    mem[16'h17C6] = 8'h06;
    mem[16'h17C7] = 8'h08;
    mem[16'h17C8] = 8'h00;
    mem[16'h17C9] = 8'h00;
    mem[16'h17CA] = 8'h00;
    mem[16'h17CB] = 8'h05; // PUSHN 8
    mem[16'h17CC] = 8'h00;
    mem[16'h17CD] = 8'h08;
    mem[16'h17CE] = 8'h00;
    mem[16'h17CF] = 8'h00;
    mem[16'h17D0] = 8'h00;
    mem[16'h17D1] = 8'h08; // POP RDI
    mem[16'h17D2] = 8'h01;
    mem[16'h17D3] = 8'h81; // ADDN RSP 8
    mem[16'h17D4] = 8'h06;
    mem[16'h17D5] = 8'h08;
    mem[16'h17D6] = 8'h00;
    mem[16'h17D7] = 8'h00;
    mem[16'h17D8] = 8'h00;
    mem[16'h17D9] = 8'h08; // POP RAX
    mem[16'h17DA] = 8'h00;
    mem[16'h17DB] = 8'h81; // ADDN RSP 8
    mem[16'h17DC] = 8'h06;
    mem[16'h17DD] = 8'h08;
    mem[16'h17DE] = 8'h00;
    mem[16'h17DF] = 8'h00;
    mem[16'h17E0] = 8'h00;
    mem[16'h17E1] = 8'h90; // CMP RAX RDI
    mem[16'h17E2] = 8'h00;
    mem[16'h17E3] = 8'h01;
    mem[16'h17E4] = 8'h18; // SETL RAX
    mem[16'h17E5] = 8'h00;
    mem[16'h17E6] = 8'h50; // MOVRR1 RAX RAX
    mem[16'h17E7] = 8'h00;
    mem[16'h17E8] = 8'h00;
    mem[16'h17E9] = 8'h85; // SUBN RSP 8
    mem[16'h17EA] = 8'h06;
    mem[16'h17EB] = 8'h08;
    mem[16'h17EC] = 8'h00;
    mem[16'h17ED] = 8'h00;
    mem[16'h17EE] = 8'h00;
    mem[16'h17EF] = 8'h04; // PUSH RAX
    mem[16'h17F0] = 8'h00;
    mem[16'h17F1] = 8'h08; // POP RAX
    mem[16'h17F2] = 8'h00;
    mem[16'h17F3] = 8'h81; // ADDN RSP 8
    mem[16'h17F4] = 8'h06;
    mem[16'h17F5] = 8'h08;
    mem[16'h17F6] = 8'h00;
    mem[16'h17F7] = 8'h00;
    mem[16'h17F8] = 8'h00;
    mem[16'h17F9] = 8'h91; // CMPN RAX 0
    mem[16'h17FA] = 8'h00;
    mem[16'h17FB] = 8'h00;
    mem[16'h17FC] = 8'h00;
    mem[16'h17FD] = 8'h00;
    mem[16'h17FE] = 8'h00;
    mem[16'h17FF] = 8'h26; // JE .Lend15
    mem[16'h1800] = 8'h16;
    mem[16'h1801] = 8'h1C;
    mem[16'h1802] = 8'h00;
    mem[16'h1803] = 8'h00;
    mem[16'h1804] = 8'h00;
    mem[16'h1805] = 8'h00;
    mem[16'h1806] = 8'h00;
    mem[16'h1807] = 8'h00;
    mem[16'h1808] = 8'h40; // MOV RAX RBP
    mem[16'h1809] = 8'h00;
    mem[16'h180A] = 8'h05;
    mem[16'h180B] = 8'h85; // SUBN RAX 8
    mem[16'h180C] = 8'h00;
    mem[16'h180D] = 8'h08;
    mem[16'h180E] = 8'h00;
    mem[16'h180F] = 8'h00;
    mem[16'h1810] = 8'h00;
    mem[16'h1811] = 8'h85; // SUBN RSP 8
    mem[16'h1812] = 8'h06;
    mem[16'h1813] = 8'h08;
    mem[16'h1814] = 8'h00;
    mem[16'h1815] = 8'h00;
    mem[16'h1816] = 8'h00;
    mem[16'h1817] = 8'h04; // PUSH RAX
    mem[16'h1818] = 8'h00;
    mem[16'h1819] = 8'h08; // POP RAX
    mem[16'h181A] = 8'h00;
    mem[16'h181B] = 8'h81; // ADDN RSP 8
    mem[16'h181C] = 8'h06;
    mem[16'h181D] = 8'h08;
    mem[16'h181E] = 8'h00;
    mem[16'h181F] = 8'h00;
    mem[16'h1820] = 8'h00;
    mem[16'h1821] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1822] = 8'h00;
    mem[16'h1823] = 8'h00;
    mem[16'h1824] = 8'h85; // SUBN RSP 8
    mem[16'h1825] = 8'h06;
    mem[16'h1826] = 8'h08;
    mem[16'h1827] = 8'h00;
    mem[16'h1828] = 8'h00;
    mem[16'h1829] = 8'h00;
    mem[16'h182A] = 8'h04; // PUSH RAX
    mem[16'h182B] = 8'h00;
    mem[16'h182C] = 8'h40; // MOV RAX RBP
    mem[16'h182D] = 8'h00;
    mem[16'h182E] = 8'h05;
    mem[16'h182F] = 8'h85; // SUBN RAX 4
    mem[16'h1830] = 8'h00;
    mem[16'h1831] = 8'h04;
    mem[16'h1832] = 8'h00;
    mem[16'h1833] = 8'h00;
    mem[16'h1834] = 8'h00;
    mem[16'h1835] = 8'h85; // SUBN RSP 8
    mem[16'h1836] = 8'h06;
    mem[16'h1837] = 8'h08;
    mem[16'h1838] = 8'h00;
    mem[16'h1839] = 8'h00;
    mem[16'h183A] = 8'h00;
    mem[16'h183B] = 8'h04; // PUSH RAX
    mem[16'h183C] = 8'h00;
    mem[16'h183D] = 8'h08; // POP RAX
    mem[16'h183E] = 8'h00;
    mem[16'h183F] = 8'h81; // ADDN RSP 8
    mem[16'h1840] = 8'h06;
    mem[16'h1841] = 8'h08;
    mem[16'h1842] = 8'h00;
    mem[16'h1843] = 8'h00;
    mem[16'h1844] = 8'h00;
    mem[16'h1845] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1846] = 8'h00;
    mem[16'h1847] = 8'h00;
    mem[16'h1848] = 8'h85; // SUBN RSP 8
    mem[16'h1849] = 8'h06;
    mem[16'h184A] = 8'h08;
    mem[16'h184B] = 8'h00;
    mem[16'h184C] = 8'h00;
    mem[16'h184D] = 8'h00;
    mem[16'h184E] = 8'h04; // PUSH RAX
    mem[16'h184F] = 8'h00;
    mem[16'h1850] = 8'h40; // MOV RAX RBP
    mem[16'h1851] = 8'h00;
    mem[16'h1852] = 8'h05;
    mem[16'h1853] = 8'h85; // SUBN RAX 12
    mem[16'h1854] = 8'h00;
    mem[16'h1855] = 8'h0C;
    mem[16'h1856] = 8'h00;
    mem[16'h1857] = 8'h00;
    mem[16'h1858] = 8'h00;
    mem[16'h1859] = 8'h85; // SUBN RSP 8
    mem[16'h185A] = 8'h06;
    mem[16'h185B] = 8'h08;
    mem[16'h185C] = 8'h00;
    mem[16'h185D] = 8'h00;
    mem[16'h185E] = 8'h00;
    mem[16'h185F] = 8'h04; // PUSH RAX
    mem[16'h1860] = 8'h00;
    mem[16'h1861] = 8'h08; // POP RAX
    mem[16'h1862] = 8'h00;
    mem[16'h1863] = 8'h81; // ADDN RSP 8
    mem[16'h1864] = 8'h06;
    mem[16'h1865] = 8'h08;
    mem[16'h1866] = 8'h00;
    mem[16'h1867] = 8'h00;
    mem[16'h1868] = 8'h00;
    mem[16'h1869] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h186A] = 8'h00;
    mem[16'h186B] = 8'h00;
    mem[16'h186C] = 8'h85; // SUBN RSP 8
    mem[16'h186D] = 8'h06;
    mem[16'h186E] = 8'h08;
    mem[16'h186F] = 8'h00;
    mem[16'h1870] = 8'h00;
    mem[16'h1871] = 8'h00;
    mem[16'h1872] = 8'h04; // PUSH RAX
    mem[16'h1873] = 8'h00;
    mem[16'h1874] = 8'h08; // POP RDX
    mem[16'h1875] = 8'h03;
    mem[16'h1876] = 8'h81; // ADDN RSP 8
    mem[16'h1877] = 8'h06;
    mem[16'h1878] = 8'h08;
    mem[16'h1879] = 8'h00;
    mem[16'h187A] = 8'h00;
    mem[16'h187B] = 8'h00;
    mem[16'h187C] = 8'h08; // POP RSI
    mem[16'h187D] = 8'h02;
    mem[16'h187E] = 8'h81; // ADDN RSP 8
    mem[16'h187F] = 8'h06;
    mem[16'h1880] = 8'h08;
    mem[16'h1881] = 8'h00;
    mem[16'h1882] = 8'h00;
    mem[16'h1883] = 8'h00;
    mem[16'h1884] = 8'h08; // POP RDI
    mem[16'h1885] = 8'h01;
    mem[16'h1886] = 8'h81; // ADDN RSP 8
    mem[16'h1887] = 8'h06;
    mem[16'h1888] = 8'h08;
    mem[16'h1889] = 8'h00;
    mem[16'h188A] = 8'h00;
    mem[16'h188B] = 8'h00;
    mem[16'h188C] = 8'h40; // MOV RAX RSP
    mem[16'h188D] = 8'h00;
    mem[16'h188E] = 8'h06;
    mem[16'h188F] = 8'h8D; // ANDN RAX 15
    mem[16'h1890] = 8'h00;
    mem[16'h1891] = 8'h0F;
    mem[16'h1892] = 8'h00;
    mem[16'h1893] = 8'h00;
    mem[16'h1894] = 8'h00;
    mem[16'h1895] = 8'h2A; // JNZ .Lcall17
    mem[16'h1896] = 8'hC6;
    mem[16'h1897] = 8'h18;
    mem[16'h1898] = 8'h00;
    mem[16'h1899] = 8'h00;
    mem[16'h189A] = 8'h00;
    mem[16'h189B] = 8'h00;
    mem[16'h189C] = 8'h00;
    mem[16'h189D] = 8'h00;
    mem[16'h189E] = 8'h41; // MOVRN RAX 0
    mem[16'h189F] = 8'h00;
    mem[16'h18A0] = 8'h00;
    mem[16'h18A1] = 8'h00;
    mem[16'h18A2] = 8'h00;
    mem[16'h18A3] = 8'h00;
    mem[16'h18A4] = 8'h0C; // MOVPC RBX
    mem[16'h18A5] = 8'h07;
    mem[16'h18A6] = 8'h81; // ADDN RBX 23
    mem[16'h18A7] = 8'h07;
    mem[16'h18A8] = 8'h17;
    mem[16'h18A9] = 8'h00;
    mem[16'h18AA] = 8'h00;
    mem[16'h18AB] = 8'h00;
    mem[16'h18AC] = 8'h85; // SUBN RSP 8
    mem[16'h18AD] = 8'h06;
    mem[16'h18AE] = 8'h08;
    mem[16'h18AF] = 8'h00;
    mem[16'h18B0] = 8'h00;
    mem[16'h18B1] = 8'h00;
    mem[16'h18B2] = 8'h04; // PUSH RBX
    mem[16'h18B3] = 8'h07;
    mem[16'h18B4] = 8'h22; // JMP check
    mem[16'h18B5] = 8'h49;
    mem[16'h18B6] = 8'h00;
    mem[16'h18B7] = 8'h00;
    mem[16'h18B8] = 8'h00;
    mem[16'h18B9] = 8'h00;
    mem[16'h18BA] = 8'h00;
    mem[16'h18BB] = 8'h00;
    mem[16'h18BC] = 8'h00;
    mem[16'h18BD] = 8'h22; // JMP .Lend17
    mem[16'h18BE] = 8'hF1;
    mem[16'h18BF] = 8'h18;
    mem[16'h18C0] = 8'h00;
    mem[16'h18C1] = 8'h00;
    mem[16'h18C2] = 8'h00;
    mem[16'h18C3] = 8'h00;
    mem[16'h18C4] = 8'h00;
    mem[16'h18C5] = 8'h00;
                          // .Lcall17:
    mem[16'h18C6] = 8'h85; // SUBN RSP 8
    mem[16'h18C7] = 8'h06;
    mem[16'h18C8] = 8'h08;
    mem[16'h18C9] = 8'h00;
    mem[16'h18CA] = 8'h00;
    mem[16'h18CB] = 8'h00;
    mem[16'h18CC] = 8'h41; // MOVRN RAX 0
    mem[16'h18CD] = 8'h00;
    mem[16'h18CE] = 8'h00;
    mem[16'h18CF] = 8'h00;
    mem[16'h18D0] = 8'h00;
    mem[16'h18D1] = 8'h00;
    mem[16'h18D2] = 8'h0C; // MOVPC RBX
    mem[16'h18D3] = 8'h07;
    mem[16'h18D4] = 8'h81; // ADDN RBX 23
    mem[16'h18D5] = 8'h07;
    mem[16'h18D6] = 8'h17;
    mem[16'h18D7] = 8'h00;
    mem[16'h18D8] = 8'h00;
    mem[16'h18D9] = 8'h00;
    mem[16'h18DA] = 8'h85; // SUBN RSP 8
    mem[16'h18DB] = 8'h06;
    mem[16'h18DC] = 8'h08;
    mem[16'h18DD] = 8'h00;
    mem[16'h18DE] = 8'h00;
    mem[16'h18DF] = 8'h00;
    mem[16'h18E0] = 8'h04; // PUSH RBX
    mem[16'h18E1] = 8'h07;
    mem[16'h18E2] = 8'h22; // JMP check
    mem[16'h18E3] = 8'h49;
    mem[16'h18E4] = 8'h00;
    mem[16'h18E5] = 8'h00;
    mem[16'h18E6] = 8'h00;
    mem[16'h18E7] = 8'h00;
    mem[16'h18E8] = 8'h00;
    mem[16'h18E9] = 8'h00;
    mem[16'h18EA] = 8'h00;
    mem[16'h18EB] = 8'h81; // ADDN RSP 8
    mem[16'h18EC] = 8'h06;
    mem[16'h18ED] = 8'h08;
    mem[16'h18EE] = 8'h00;
    mem[16'h18EF] = 8'h00;
    mem[16'h18F0] = 8'h00;
                          // .Lend17:
    mem[16'h18F1] = 8'h85; // SUBN RSP 8
    mem[16'h18F2] = 8'h06;
    mem[16'h18F3] = 8'h08;
    mem[16'h18F4] = 8'h00;
    mem[16'h18F5] = 8'h00;
    mem[16'h18F6] = 8'h00;
    mem[16'h18F7] = 8'h04; // PUSH RAX
    mem[16'h18F8] = 8'h00;
    mem[16'h18F9] = 8'h08; // POP RAX
    mem[16'h18FA] = 8'h00;
    mem[16'h18FB] = 8'h81; // ADDN RSP 8
    mem[16'h18FC] = 8'h06;
    mem[16'h18FD] = 8'h08;
    mem[16'h18FE] = 8'h00;
    mem[16'h18FF] = 8'h00;
    mem[16'h1900] = 8'h00;
    mem[16'h1901] = 8'h91; // CMPN RAX 0
    mem[16'h1902] = 8'h00;
    mem[16'h1903] = 8'h00;
    mem[16'h1904] = 8'h00;
    mem[16'h1905] = 8'h00;
    mem[16'h1906] = 8'h00;
    mem[16'h1907] = 8'h26; // JE .Lend16
    mem[16'h1908] = 8'h90;
    mem[16'h1909] = 8'h1B;
    mem[16'h190A] = 8'h00;
    mem[16'h190B] = 8'h00;
    mem[16'h190C] = 8'h00;
    mem[16'h190D] = 8'h00;
    mem[16'h190E] = 8'h00;
    mem[16'h190F] = 8'h00;
    mem[16'h1910] = 8'h85; // SUBN RSP 8
    mem[16'h1911] = 8'h06;
    mem[16'h1912] = 8'h08;
    mem[16'h1913] = 8'h00;
    mem[16'h1914] = 8'h00;
    mem[16'h1915] = 8'h00;
    mem[16'h1916] = 8'h06; // PUSHA pos
    mem[16'h1917] = 8'h09;
    mem[16'h1918] = 8'h00;
    mem[16'h1919] = 8'h00;
    mem[16'h191A] = 8'h00;
    mem[16'h191B] = 8'h00;
    mem[16'h191C] = 8'h00;
    mem[16'h191D] = 8'h00;
    mem[16'h191E] = 8'h00;
    mem[16'h191F] = 8'h40; // MOV RAX RBP
    mem[16'h1920] = 8'h00;
    mem[16'h1921] = 8'h05;
    mem[16'h1922] = 8'h85; // SUBN RAX 12
    mem[16'h1923] = 8'h00;
    mem[16'h1924] = 8'h0C;
    mem[16'h1925] = 8'h00;
    mem[16'h1926] = 8'h00;
    mem[16'h1927] = 8'h00;
    mem[16'h1928] = 8'h85; // SUBN RSP 8
    mem[16'h1929] = 8'h06;
    mem[16'h192A] = 8'h08;
    mem[16'h192B] = 8'h00;
    mem[16'h192C] = 8'h00;
    mem[16'h192D] = 8'h00;
    mem[16'h192E] = 8'h04; // PUSH RAX
    mem[16'h192F] = 8'h00;
    mem[16'h1930] = 8'h08; // POP RAX
    mem[16'h1931] = 8'h00;
    mem[16'h1932] = 8'h81; // ADDN RSP 8
    mem[16'h1933] = 8'h06;
    mem[16'h1934] = 8'h08;
    mem[16'h1935] = 8'h00;
    mem[16'h1936] = 8'h00;
    mem[16'h1937] = 8'h00;
    mem[16'h1938] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1939] = 8'h00;
    mem[16'h193A] = 8'h00;
    mem[16'h193B] = 8'h85; // SUBN RSP 8
    mem[16'h193C] = 8'h06;
    mem[16'h193D] = 8'h08;
    mem[16'h193E] = 8'h00;
    mem[16'h193F] = 8'h00;
    mem[16'h1940] = 8'h00;
    mem[16'h1941] = 8'h04; // PUSH RAX
    mem[16'h1942] = 8'h00;
    mem[16'h1943] = 8'h08; // POP RDI
    mem[16'h1944] = 8'h01;
    mem[16'h1945] = 8'h81; // ADDN RSP 8
    mem[16'h1946] = 8'h06;
    mem[16'h1947] = 8'h08;
    mem[16'h1948] = 8'h00;
    mem[16'h1949] = 8'h00;
    mem[16'h194A] = 8'h00;
    mem[16'h194B] = 8'h08; // POP RAX
    mem[16'h194C] = 8'h00;
    mem[16'h194D] = 8'h81; // ADDN RSP 8
    mem[16'h194E] = 8'h06;
    mem[16'h194F] = 8'h08;
    mem[16'h1950] = 8'h00;
    mem[16'h1951] = 8'h00;
    mem[16'h1952] = 8'h00;
    mem[16'h1953] = 8'h89; // MULN RDI 8
    mem[16'h1954] = 8'h01;
    mem[16'h1955] = 8'h08;
    mem[16'h1956] = 8'h00;
    mem[16'h1957] = 8'h00;
    mem[16'h1958] = 8'h00;
    mem[16'h1959] = 8'h80; // ADD RAX RDI
    mem[16'h195A] = 8'h00;
    mem[16'h195B] = 8'h01;
    mem[16'h195C] = 8'h85; // SUBN RSP 8
    mem[16'h195D] = 8'h06;
    mem[16'h195E] = 8'h08;
    mem[16'h195F] = 8'h00;
    mem[16'h1960] = 8'h00;
    mem[16'h1961] = 8'h00;
    mem[16'h1962] = 8'h04; // PUSH RAX
    mem[16'h1963] = 8'h00;
    mem[16'h1964] = 8'h85; // SUBN RSP 8
    mem[16'h1965] = 8'h06;
    mem[16'h1966] = 8'h08;
    mem[16'h1967] = 8'h00;
    mem[16'h1968] = 8'h00;
    mem[16'h1969] = 8'h00;
    mem[16'h196A] = 8'h05; // PUSHN 0
    mem[16'h196B] = 8'h00;
    mem[16'h196C] = 8'h00;
    mem[16'h196D] = 8'h00;
    mem[16'h196E] = 8'h00;
    mem[16'h196F] = 8'h00;
    mem[16'h1970] = 8'h08; // POP RDI
    mem[16'h1971] = 8'h01;
    mem[16'h1972] = 8'h81; // ADDN RSP 8
    mem[16'h1973] = 8'h06;
    mem[16'h1974] = 8'h08;
    mem[16'h1975] = 8'h00;
    mem[16'h1976] = 8'h00;
    mem[16'h1977] = 8'h00;
    mem[16'h1978] = 8'h08; // POP RAX
    mem[16'h1979] = 8'h00;
    mem[16'h197A] = 8'h81; // ADDN RSP 8
    mem[16'h197B] = 8'h06;
    mem[16'h197C] = 8'h08;
    mem[16'h197D] = 8'h00;
    mem[16'h197E] = 8'h00;
    mem[16'h197F] = 8'h00;
    mem[16'h1980] = 8'h89; // MULN RDI 4
    mem[16'h1981] = 8'h01;
    mem[16'h1982] = 8'h04;
    mem[16'h1983] = 8'h00;
    mem[16'h1984] = 8'h00;
    mem[16'h1985] = 8'h00;
    mem[16'h1986] = 8'h80; // ADD RAX RDI
    mem[16'h1987] = 8'h00;
    mem[16'h1988] = 8'h01;
    mem[16'h1989] = 8'h85; // SUBN RSP 8
    mem[16'h198A] = 8'h06;
    mem[16'h198B] = 8'h08;
    mem[16'h198C] = 8'h00;
    mem[16'h198D] = 8'h00;
    mem[16'h198E] = 8'h00;
    mem[16'h198F] = 8'h04; // PUSH RAX
    mem[16'h1990] = 8'h00;
    mem[16'h1991] = 8'h40; // MOV RAX RBP
    mem[16'h1992] = 8'h00;
    mem[16'h1993] = 8'h05;
    mem[16'h1994] = 8'h85; // SUBN RAX 8
    mem[16'h1995] = 8'h00;
    mem[16'h1996] = 8'h08;
    mem[16'h1997] = 8'h00;
    mem[16'h1998] = 8'h00;
    mem[16'h1999] = 8'h00;
    mem[16'h199A] = 8'h85; // SUBN RSP 8
    mem[16'h199B] = 8'h06;
    mem[16'h199C] = 8'h08;
    mem[16'h199D] = 8'h00;
    mem[16'h199E] = 8'h00;
    mem[16'h199F] = 8'h00;
    mem[16'h19A0] = 8'h04; // PUSH RAX
    mem[16'h19A1] = 8'h00;
    mem[16'h19A2] = 8'h08; // POP RAX
    mem[16'h19A3] = 8'h00;
    mem[16'h19A4] = 8'h81; // ADDN RSP 8
    mem[16'h19A5] = 8'h06;
    mem[16'h19A6] = 8'h08;
    mem[16'h19A7] = 8'h00;
    mem[16'h19A8] = 8'h00;
    mem[16'h19A9] = 8'h00;
    mem[16'h19AA] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h19AB] = 8'h00;
    mem[16'h19AC] = 8'h00;
    mem[16'h19AD] = 8'h85; // SUBN RSP 8
    mem[16'h19AE] = 8'h06;
    mem[16'h19AF] = 8'h08;
    mem[16'h19B0] = 8'h00;
    mem[16'h19B1] = 8'h00;
    mem[16'h19B2] = 8'h00;
    mem[16'h19B3] = 8'h04; // PUSH RAX
    mem[16'h19B4] = 8'h00;
    mem[16'h19B5] = 8'h08; // POP RDI
    mem[16'h19B6] = 8'h01;
    mem[16'h19B7] = 8'h81; // ADDN RSP 8
    mem[16'h19B8] = 8'h06;
    mem[16'h19B9] = 8'h08;
    mem[16'h19BA] = 8'h00;
    mem[16'h19BB] = 8'h00;
    mem[16'h19BC] = 8'h00;
    mem[16'h19BD] = 8'h08; // POP RAX
    mem[16'h19BE] = 8'h00;
    mem[16'h19BF] = 8'h81; // ADDN RSP 8
    mem[16'h19C0] = 8'h06;
    mem[16'h19C1] = 8'h08;
    mem[16'h19C2] = 8'h00;
    mem[16'h19C3] = 8'h00;
    mem[16'h19C4] = 8'h00;
    mem[16'h19C5] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h19C6] = 8'h00;
    mem[16'h19C7] = 8'h01;
    mem[16'h19C8] = 8'h85; // SUBN RSP 8
    mem[16'h19C9] = 8'h06;
    mem[16'h19CA] = 8'h08;
    mem[16'h19CB] = 8'h00;
    mem[16'h19CC] = 8'h00;
    mem[16'h19CD] = 8'h00;
    mem[16'h19CE] = 8'h04; // PUSH RDI
    mem[16'h19CF] = 8'h01;
    mem[16'h19D0] = 8'h81; // ADDN RSP 8
    mem[16'h19D1] = 8'h06;
    mem[16'h19D2] = 8'h08;
    mem[16'h19D3] = 8'h00;
    mem[16'h19D4] = 8'h00;
    mem[16'h19D5] = 8'h00;
    mem[16'h19D6] = 8'h85; // SUBN RSP 8
    mem[16'h19D7] = 8'h06;
    mem[16'h19D8] = 8'h08;
    mem[16'h19D9] = 8'h00;
    mem[16'h19DA] = 8'h00;
    mem[16'h19DB] = 8'h00;
    mem[16'h19DC] = 8'h06; // PUSHA pos
    mem[16'h19DD] = 8'h09;
    mem[16'h19DE] = 8'h00;
    mem[16'h19DF] = 8'h00;
    mem[16'h19E0] = 8'h00;
    mem[16'h19E1] = 8'h00;
    mem[16'h19E2] = 8'h00;
    mem[16'h19E3] = 8'h00;
    mem[16'h19E4] = 8'h00;
    mem[16'h19E5] = 8'h40; // MOV RAX RBP
    mem[16'h19E6] = 8'h00;
    mem[16'h19E7] = 8'h05;
    mem[16'h19E8] = 8'h85; // SUBN RAX 12
    mem[16'h19E9] = 8'h00;
    mem[16'h19EA] = 8'h0C;
    mem[16'h19EB] = 8'h00;
    mem[16'h19EC] = 8'h00;
    mem[16'h19ED] = 8'h00;
    mem[16'h19EE] = 8'h85; // SUBN RSP 8
    mem[16'h19EF] = 8'h06;
    mem[16'h19F0] = 8'h08;
    mem[16'h19F1] = 8'h00;
    mem[16'h19F2] = 8'h00;
    mem[16'h19F3] = 8'h00;
    mem[16'h19F4] = 8'h04; // PUSH RAX
    mem[16'h19F5] = 8'h00;
    mem[16'h19F6] = 8'h08; // POP RAX
    mem[16'h19F7] = 8'h00;
    mem[16'h19F8] = 8'h81; // ADDN RSP 8
    mem[16'h19F9] = 8'h06;
    mem[16'h19FA] = 8'h08;
    mem[16'h19FB] = 8'h00;
    mem[16'h19FC] = 8'h00;
    mem[16'h19FD] = 8'h00;
    mem[16'h19FE] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h19FF] = 8'h00;
    mem[16'h1A00] = 8'h00;
    mem[16'h1A01] = 8'h85; // SUBN RSP 8
    mem[16'h1A02] = 8'h06;
    mem[16'h1A03] = 8'h08;
    mem[16'h1A04] = 8'h00;
    mem[16'h1A05] = 8'h00;
    mem[16'h1A06] = 8'h00;
    mem[16'h1A07] = 8'h04; // PUSH RAX
    mem[16'h1A08] = 8'h00;
    mem[16'h1A09] = 8'h08; // POP RDI
    mem[16'h1A0A] = 8'h01;
    mem[16'h1A0B] = 8'h81; // ADDN RSP 8
    mem[16'h1A0C] = 8'h06;
    mem[16'h1A0D] = 8'h08;
    mem[16'h1A0E] = 8'h00;
    mem[16'h1A0F] = 8'h00;
    mem[16'h1A10] = 8'h00;
    mem[16'h1A11] = 8'h08; // POP RAX
    mem[16'h1A12] = 8'h00;
    mem[16'h1A13] = 8'h81; // ADDN RSP 8
    mem[16'h1A14] = 8'h06;
    mem[16'h1A15] = 8'h08;
    mem[16'h1A16] = 8'h00;
    mem[16'h1A17] = 8'h00;
    mem[16'h1A18] = 8'h00;
    mem[16'h1A19] = 8'h89; // MULN RDI 8
    mem[16'h1A1A] = 8'h01;
    mem[16'h1A1B] = 8'h08;
    mem[16'h1A1C] = 8'h00;
    mem[16'h1A1D] = 8'h00;
    mem[16'h1A1E] = 8'h00;
    mem[16'h1A1F] = 8'h80; // ADD RAX RDI
    mem[16'h1A20] = 8'h00;
    mem[16'h1A21] = 8'h01;
    mem[16'h1A22] = 8'h85; // SUBN RSP 8
    mem[16'h1A23] = 8'h06;
    mem[16'h1A24] = 8'h08;
    mem[16'h1A25] = 8'h00;
    mem[16'h1A26] = 8'h00;
    mem[16'h1A27] = 8'h00;
    mem[16'h1A28] = 8'h04; // PUSH RAX
    mem[16'h1A29] = 8'h00;
    mem[16'h1A2A] = 8'h85; // SUBN RSP 8
    mem[16'h1A2B] = 8'h06;
    mem[16'h1A2C] = 8'h08;
    mem[16'h1A2D] = 8'h00;
    mem[16'h1A2E] = 8'h00;
    mem[16'h1A2F] = 8'h00;
    mem[16'h1A30] = 8'h05; // PUSHN 1
    mem[16'h1A31] = 8'h00;
    mem[16'h1A32] = 8'h01;
    mem[16'h1A33] = 8'h00;
    mem[16'h1A34] = 8'h00;
    mem[16'h1A35] = 8'h00;
    mem[16'h1A36] = 8'h08; // POP RDI
    mem[16'h1A37] = 8'h01;
    mem[16'h1A38] = 8'h81; // ADDN RSP 8
    mem[16'h1A39] = 8'h06;
    mem[16'h1A3A] = 8'h08;
    mem[16'h1A3B] = 8'h00;
    mem[16'h1A3C] = 8'h00;
    mem[16'h1A3D] = 8'h00;
    mem[16'h1A3E] = 8'h08; // POP RAX
    mem[16'h1A3F] = 8'h00;
    mem[16'h1A40] = 8'h81; // ADDN RSP 8
    mem[16'h1A41] = 8'h06;
    mem[16'h1A42] = 8'h08;
    mem[16'h1A43] = 8'h00;
    mem[16'h1A44] = 8'h00;
    mem[16'h1A45] = 8'h00;
    mem[16'h1A46] = 8'h89; // MULN RDI 4
    mem[16'h1A47] = 8'h01;
    mem[16'h1A48] = 8'h04;
    mem[16'h1A49] = 8'h00;
    mem[16'h1A4A] = 8'h00;
    mem[16'h1A4B] = 8'h00;
    mem[16'h1A4C] = 8'h80; // ADD RAX RDI
    mem[16'h1A4D] = 8'h00;
    mem[16'h1A4E] = 8'h01;
    mem[16'h1A4F] = 8'h85; // SUBN RSP 8
    mem[16'h1A50] = 8'h06;
    mem[16'h1A51] = 8'h08;
    mem[16'h1A52] = 8'h00;
    mem[16'h1A53] = 8'h00;
    mem[16'h1A54] = 8'h00;
    mem[16'h1A55] = 8'h04; // PUSH RAX
    mem[16'h1A56] = 8'h00;
    mem[16'h1A57] = 8'h40; // MOV RAX RBP
    mem[16'h1A58] = 8'h00;
    mem[16'h1A59] = 8'h05;
    mem[16'h1A5A] = 8'h85; // SUBN RAX 4
    mem[16'h1A5B] = 8'h00;
    mem[16'h1A5C] = 8'h04;
    mem[16'h1A5D] = 8'h00;
    mem[16'h1A5E] = 8'h00;
    mem[16'h1A5F] = 8'h00;
    mem[16'h1A60] = 8'h85; // SUBN RSP 8
    mem[16'h1A61] = 8'h06;
    mem[16'h1A62] = 8'h08;
    mem[16'h1A63] = 8'h00;
    mem[16'h1A64] = 8'h00;
    mem[16'h1A65] = 8'h00;
    mem[16'h1A66] = 8'h04; // PUSH RAX
    mem[16'h1A67] = 8'h00;
    mem[16'h1A68] = 8'h08; // POP RAX
    mem[16'h1A69] = 8'h00;
    mem[16'h1A6A] = 8'h81; // ADDN RSP 8
    mem[16'h1A6B] = 8'h06;
    mem[16'h1A6C] = 8'h08;
    mem[16'h1A6D] = 8'h00;
    mem[16'h1A6E] = 8'h00;
    mem[16'h1A6F] = 8'h00;
    mem[16'h1A70] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1A71] = 8'h00;
    mem[16'h1A72] = 8'h00;
    mem[16'h1A73] = 8'h85; // SUBN RSP 8
    mem[16'h1A74] = 8'h06;
    mem[16'h1A75] = 8'h08;
    mem[16'h1A76] = 8'h00;
    mem[16'h1A77] = 8'h00;
    mem[16'h1A78] = 8'h00;
    mem[16'h1A79] = 8'h04; // PUSH RAX
    mem[16'h1A7A] = 8'h00;
    mem[16'h1A7B] = 8'h08; // POP RDI
    mem[16'h1A7C] = 8'h01;
    mem[16'h1A7D] = 8'h81; // ADDN RSP 8
    mem[16'h1A7E] = 8'h06;
    mem[16'h1A7F] = 8'h08;
    mem[16'h1A80] = 8'h00;
    mem[16'h1A81] = 8'h00;
    mem[16'h1A82] = 8'h00;
    mem[16'h1A83] = 8'h08; // POP RAX
    mem[16'h1A84] = 8'h00;
    mem[16'h1A85] = 8'h81; // ADDN RSP 8
    mem[16'h1A86] = 8'h06;
    mem[16'h1A87] = 8'h08;
    mem[16'h1A88] = 8'h00;
    mem[16'h1A89] = 8'h00;
    mem[16'h1A8A] = 8'h00;
    mem[16'h1A8B] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h1A8C] = 8'h00;
    mem[16'h1A8D] = 8'h01;
    mem[16'h1A8E] = 8'h85; // SUBN RSP 8
    mem[16'h1A8F] = 8'h06;
    mem[16'h1A90] = 8'h08;
    mem[16'h1A91] = 8'h00;
    mem[16'h1A92] = 8'h00;
    mem[16'h1A93] = 8'h00;
    mem[16'h1A94] = 8'h04; // PUSH RDI
    mem[16'h1A95] = 8'h01;
    mem[16'h1A96] = 8'h81; // ADDN RSP 8
    mem[16'h1A97] = 8'h06;
    mem[16'h1A98] = 8'h08;
    mem[16'h1A99] = 8'h00;
    mem[16'h1A9A] = 8'h00;
    mem[16'h1A9B] = 8'h00;
    mem[16'h1A9C] = 8'h40; // MOV RAX RBP
    mem[16'h1A9D] = 8'h00;
    mem[16'h1A9E] = 8'h05;
    mem[16'h1A9F] = 8'h85; // SUBN RAX 12
    mem[16'h1AA0] = 8'h00;
    mem[16'h1AA1] = 8'h0C;
    mem[16'h1AA2] = 8'h00;
    mem[16'h1AA3] = 8'h00;
    mem[16'h1AA4] = 8'h00;
    mem[16'h1AA5] = 8'h85; // SUBN RSP 8
    mem[16'h1AA6] = 8'h06;
    mem[16'h1AA7] = 8'h08;
    mem[16'h1AA8] = 8'h00;
    mem[16'h1AA9] = 8'h00;
    mem[16'h1AAA] = 8'h00;
    mem[16'h1AAB] = 8'h04; // PUSH RAX
    mem[16'h1AAC] = 8'h00;
    mem[16'h1AAD] = 8'h08; // POP RAX
    mem[16'h1AAE] = 8'h00;
    mem[16'h1AAF] = 8'h81; // ADDN RSP 8
    mem[16'h1AB0] = 8'h06;
    mem[16'h1AB1] = 8'h08;
    mem[16'h1AB2] = 8'h00;
    mem[16'h1AB3] = 8'h00;
    mem[16'h1AB4] = 8'h00;
    mem[16'h1AB5] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1AB6] = 8'h00;
    mem[16'h1AB7] = 8'h00;
    mem[16'h1AB8] = 8'h85; // SUBN RSP 8
    mem[16'h1AB9] = 8'h06;
    mem[16'h1ABA] = 8'h08;
    mem[16'h1ABB] = 8'h00;
    mem[16'h1ABC] = 8'h00;
    mem[16'h1ABD] = 8'h00;
    mem[16'h1ABE] = 8'h04; // PUSH RAX
    mem[16'h1ABF] = 8'h00;
    mem[16'h1AC0] = 8'h85; // SUBN RSP 8
    mem[16'h1AC1] = 8'h06;
    mem[16'h1AC2] = 8'h08;
    mem[16'h1AC3] = 8'h00;
    mem[16'h1AC4] = 8'h00;
    mem[16'h1AC5] = 8'h00;
    mem[16'h1AC6] = 8'h05; // PUSHN 1
    mem[16'h1AC7] = 8'h00;
    mem[16'h1AC8] = 8'h01;
    mem[16'h1AC9] = 8'h00;
    mem[16'h1ACA] = 8'h00;
    mem[16'h1ACB] = 8'h00;
    mem[16'h1ACC] = 8'h08; // POP RDI
    mem[16'h1ACD] = 8'h01;
    mem[16'h1ACE] = 8'h81; // ADDN RSP 8
    mem[16'h1ACF] = 8'h06;
    mem[16'h1AD0] = 8'h08;
    mem[16'h1AD1] = 8'h00;
    mem[16'h1AD2] = 8'h00;
    mem[16'h1AD3] = 8'h00;
    mem[16'h1AD4] = 8'h08; // POP RAX
    mem[16'h1AD5] = 8'h00;
    mem[16'h1AD6] = 8'h81; // ADDN RSP 8
    mem[16'h1AD7] = 8'h06;
    mem[16'h1AD8] = 8'h08;
    mem[16'h1AD9] = 8'h00;
    mem[16'h1ADA] = 8'h00;
    mem[16'h1ADB] = 8'h00;
    mem[16'h1ADC] = 8'h80; // ADD RAX RDI
    mem[16'h1ADD] = 8'h00;
    mem[16'h1ADE] = 8'h01;
    mem[16'h1ADF] = 8'h85; // SUBN RSP 8
    mem[16'h1AE0] = 8'h06;
    mem[16'h1AE1] = 8'h08;
    mem[16'h1AE2] = 8'h00;
    mem[16'h1AE3] = 8'h00;
    mem[16'h1AE4] = 8'h00;
    mem[16'h1AE5] = 8'h04; // PUSH RAX
    mem[16'h1AE6] = 8'h00;
    mem[16'h1AE7] = 8'h08; // POP RDI
    mem[16'h1AE8] = 8'h01;
    mem[16'h1AE9] = 8'h81; // ADDN RSP 8
    mem[16'h1AEA] = 8'h06;
    mem[16'h1AEB] = 8'h08;
    mem[16'h1AEC] = 8'h00;
    mem[16'h1AED] = 8'h00;
    mem[16'h1AEE] = 8'h00;
    mem[16'h1AEF] = 8'h40; // MOV RAX RSP
    mem[16'h1AF0] = 8'h00;
    mem[16'h1AF1] = 8'h06;
    mem[16'h1AF2] = 8'h8D; // ANDN RAX 15
    mem[16'h1AF3] = 8'h00;
    mem[16'h1AF4] = 8'h0F;
    mem[16'h1AF5] = 8'h00;
    mem[16'h1AF6] = 8'h00;
    mem[16'h1AF7] = 8'h00;
    mem[16'h1AF8] = 8'h2A; // JNZ .Lcall19
    mem[16'h1AF9] = 8'h29;
    mem[16'h1AFA] = 8'h1B;
    mem[16'h1AFB] = 8'h00;
    mem[16'h1AFC] = 8'h00;
    mem[16'h1AFD] = 8'h00;
    mem[16'h1AFE] = 8'h00;
    mem[16'h1AFF] = 8'h00;
    mem[16'h1B00] = 8'h00;
    mem[16'h1B01] = 8'h41; // MOVRN RAX 0
    mem[16'h1B02] = 8'h00;
    mem[16'h1B03] = 8'h00;
    mem[16'h1B04] = 8'h00;
    mem[16'h1B05] = 8'h00;
    mem[16'h1B06] = 8'h00;
    mem[16'h1B07] = 8'h0C; // MOVPC RBX
    mem[16'h1B08] = 8'h07;
    mem[16'h1B09] = 8'h81; // ADDN RBX 23
    mem[16'h1B0A] = 8'h07;
    mem[16'h1B0B] = 8'h17;
    mem[16'h1B0C] = 8'h00;
    mem[16'h1B0D] = 8'h00;
    mem[16'h1B0E] = 8'h00;
    mem[16'h1B0F] = 8'h85; // SUBN RSP 8
    mem[16'h1B10] = 8'h06;
    mem[16'h1B11] = 8'h08;
    mem[16'h1B12] = 8'h00;
    mem[16'h1B13] = 8'h00;
    mem[16'h1B14] = 8'h00;
    mem[16'h1B15] = 8'h04; // PUSH RBX
    mem[16'h1B16] = 8'h07;
    mem[16'h1B17] = 8'h22; // JMP eightqueen
    mem[16'h1B18] = 8'h1D;
    mem[16'h1B19] = 8'h16;
    mem[16'h1B1A] = 8'h00;
    mem[16'h1B1B] = 8'h00;
    mem[16'h1B1C] = 8'h00;
    mem[16'h1B1D] = 8'h00;
    mem[16'h1B1E] = 8'h00;
    mem[16'h1B1F] = 8'h00;
    mem[16'h1B20] = 8'h22; // JMP .Lend19
    mem[16'h1B21] = 8'h54;
    mem[16'h1B22] = 8'h1B;
    mem[16'h1B23] = 8'h00;
    mem[16'h1B24] = 8'h00;
    mem[16'h1B25] = 8'h00;
    mem[16'h1B26] = 8'h00;
    mem[16'h1B27] = 8'h00;
    mem[16'h1B28] = 8'h00;
                          // .Lcall19:
    mem[16'h1B29] = 8'h85; // SUBN RSP 8
    mem[16'h1B2A] = 8'h06;
    mem[16'h1B2B] = 8'h08;
    mem[16'h1B2C] = 8'h00;
    mem[16'h1B2D] = 8'h00;
    mem[16'h1B2E] = 8'h00;
    mem[16'h1B2F] = 8'h41; // MOVRN RAX 0
    mem[16'h1B30] = 8'h00;
    mem[16'h1B31] = 8'h00;
    mem[16'h1B32] = 8'h00;
    mem[16'h1B33] = 8'h00;
    mem[16'h1B34] = 8'h00;
    mem[16'h1B35] = 8'h0C; // MOVPC RBX
    mem[16'h1B36] = 8'h07;
    mem[16'h1B37] = 8'h81; // ADDN RBX 23
    mem[16'h1B38] = 8'h07;
    mem[16'h1B39] = 8'h17;
    mem[16'h1B3A] = 8'h00;
    mem[16'h1B3B] = 8'h00;
    mem[16'h1B3C] = 8'h00;
    mem[16'h1B3D] = 8'h85; // SUBN RSP 8
    mem[16'h1B3E] = 8'h06;
    mem[16'h1B3F] = 8'h08;
    mem[16'h1B40] = 8'h00;
    mem[16'h1B41] = 8'h00;
    mem[16'h1B42] = 8'h00;
    mem[16'h1B43] = 8'h04; // PUSH RBX
    mem[16'h1B44] = 8'h07;
    mem[16'h1B45] = 8'h22; // JMP eightqueen
    mem[16'h1B46] = 8'h1D;
    mem[16'h1B47] = 8'h16;
    mem[16'h1B48] = 8'h00;
    mem[16'h1B49] = 8'h00;
    mem[16'h1B4A] = 8'h00;
    mem[16'h1B4B] = 8'h00;
    mem[16'h1B4C] = 8'h00;
    mem[16'h1B4D] = 8'h00;
    mem[16'h1B4E] = 8'h81; // ADDN RSP 8
    mem[16'h1B4F] = 8'h06;
    mem[16'h1B50] = 8'h08;
    mem[16'h1B51] = 8'h00;
    mem[16'h1B52] = 8'h00;
    mem[16'h1B53] = 8'h00;
                          // .Lend19:
    mem[16'h1B54] = 8'h85; // SUBN RSP 8
    mem[16'h1B55] = 8'h06;
    mem[16'h1B56] = 8'h08;
    mem[16'h1B57] = 8'h00;
    mem[16'h1B58] = 8'h00;
    mem[16'h1B59] = 8'h00;
    mem[16'h1B5A] = 8'h04; // PUSH RAX
    mem[16'h1B5B] = 8'h00;
    mem[16'h1B5C] = 8'h08; // POP RAX
    mem[16'h1B5D] = 8'h00;
    mem[16'h1B5E] = 8'h81; // ADDN RSP 8
    mem[16'h1B5F] = 8'h06;
    mem[16'h1B60] = 8'h08;
    mem[16'h1B61] = 8'h00;
    mem[16'h1B62] = 8'h00;
    mem[16'h1B63] = 8'h00;
    mem[16'h1B64] = 8'h91; // CMPN RAX 0
    mem[16'h1B65] = 8'h00;
    mem[16'h1B66] = 8'h00;
    mem[16'h1B67] = 8'h00;
    mem[16'h1B68] = 8'h00;
    mem[16'h1B69] = 8'h00;
    mem[16'h1B6A] = 8'h26; // JE .Lend18
    mem[16'h1B6B] = 8'h90;
    mem[16'h1B6C] = 8'h1B;
    mem[16'h1B6D] = 8'h00;
    mem[16'h1B6E] = 8'h00;
    mem[16'h1B6F] = 8'h00;
    mem[16'h1B70] = 8'h00;
    mem[16'h1B71] = 8'h00;
    mem[16'h1B72] = 8'h00;
    mem[16'h1B73] = 8'h85; // SUBN RSP 8
    mem[16'h1B74] = 8'h06;
    mem[16'h1B75] = 8'h08;
    mem[16'h1B76] = 8'h00;
    mem[16'h1B77] = 8'h00;
    mem[16'h1B78] = 8'h00;
    mem[16'h1B79] = 8'h05; // PUSHN 1
    mem[16'h1B7A] = 8'h00;
    mem[16'h1B7B] = 8'h01;
    mem[16'h1B7C] = 8'h00;
    mem[16'h1B7D] = 8'h00;
    mem[16'h1B7E] = 8'h00;
    mem[16'h1B7F] = 8'h08; // POP RAX
    mem[16'h1B80] = 8'h00;
    mem[16'h1B81] = 8'h81; // ADDN RSP 8
    mem[16'h1B82] = 8'h06;
    mem[16'h1B83] = 8'h08;
    mem[16'h1B84] = 8'h00;
    mem[16'h1B85] = 8'h00;
    mem[16'h1B86] = 8'h00;
    mem[16'h1B87] = 8'h22; // JMP .Lreturn.eightqueen
    mem[16'h1B88] = 8'hB9;
    mem[16'h1B89] = 8'h1C;
    mem[16'h1B8A] = 8'h00;
    mem[16'h1B8B] = 8'h00;
    mem[16'h1B8C] = 8'h00;
    mem[16'h1B8D] = 8'h00;
    mem[16'h1B8E] = 8'h00;
    mem[16'h1B8F] = 8'h00;
                          // .Lend18:
                          // .Lend16:
    mem[16'h1B90] = 8'h40; // MOV RAX RBP
    mem[16'h1B91] = 8'h00;
    mem[16'h1B92] = 8'h05;
    mem[16'h1B93] = 8'h85; // SUBN RAX 8
    mem[16'h1B94] = 8'h00;
    mem[16'h1B95] = 8'h08;
    mem[16'h1B96] = 8'h00;
    mem[16'h1B97] = 8'h00;
    mem[16'h1B98] = 8'h00;
    mem[16'h1B99] = 8'h85; // SUBN RSP 8
    mem[16'h1B9A] = 8'h06;
    mem[16'h1B9B] = 8'h08;
    mem[16'h1B9C] = 8'h00;
    mem[16'h1B9D] = 8'h00;
    mem[16'h1B9E] = 8'h00;
    mem[16'h1B9F] = 8'h04; // PUSH RAX
    mem[16'h1BA0] = 8'h00;
    mem[16'h1BA1] = 8'h40; // MOV RAX RBP
    mem[16'h1BA2] = 8'h00;
    mem[16'h1BA3] = 8'h05;
    mem[16'h1BA4] = 8'h85; // SUBN RAX 8
    mem[16'h1BA5] = 8'h00;
    mem[16'h1BA6] = 8'h08;
    mem[16'h1BA7] = 8'h00;
    mem[16'h1BA8] = 8'h00;
    mem[16'h1BA9] = 8'h00;
    mem[16'h1BAA] = 8'h85; // SUBN RSP 8
    mem[16'h1BAB] = 8'h06;
    mem[16'h1BAC] = 8'h08;
    mem[16'h1BAD] = 8'h00;
    mem[16'h1BAE] = 8'h00;
    mem[16'h1BAF] = 8'h00;
    mem[16'h1BB0] = 8'h04; // PUSH RAX
    mem[16'h1BB1] = 8'h00;
    mem[16'h1BB2] = 8'h08; // POP RAX
    mem[16'h1BB3] = 8'h00;
    mem[16'h1BB4] = 8'h81; // ADDN RSP 8
    mem[16'h1BB5] = 8'h06;
    mem[16'h1BB6] = 8'h08;
    mem[16'h1BB7] = 8'h00;
    mem[16'h1BB8] = 8'h00;
    mem[16'h1BB9] = 8'h00;
    mem[16'h1BBA] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1BBB] = 8'h00;
    mem[16'h1BBC] = 8'h00;
    mem[16'h1BBD] = 8'h85; // SUBN RSP 8
    mem[16'h1BBE] = 8'h06;
    mem[16'h1BBF] = 8'h08;
    mem[16'h1BC0] = 8'h00;
    mem[16'h1BC1] = 8'h00;
    mem[16'h1BC2] = 8'h00;
    mem[16'h1BC3] = 8'h04; // PUSH RAX
    mem[16'h1BC4] = 8'h00;
    mem[16'h1BC5] = 8'h85; // SUBN RSP 8
    mem[16'h1BC6] = 8'h06;
    mem[16'h1BC7] = 8'h08;
    mem[16'h1BC8] = 8'h00;
    mem[16'h1BC9] = 8'h00;
    mem[16'h1BCA] = 8'h00;
    mem[16'h1BCB] = 8'h05; // PUSHN 1
    mem[16'h1BCC] = 8'h00;
    mem[16'h1BCD] = 8'h01;
    mem[16'h1BCE] = 8'h00;
    mem[16'h1BCF] = 8'h00;
    mem[16'h1BD0] = 8'h00;
    mem[16'h1BD1] = 8'h08; // POP RDI
    mem[16'h1BD2] = 8'h01;
    mem[16'h1BD3] = 8'h81; // ADDN RSP 8
    mem[16'h1BD4] = 8'h06;
    mem[16'h1BD5] = 8'h08;
    mem[16'h1BD6] = 8'h00;
    mem[16'h1BD7] = 8'h00;
    mem[16'h1BD8] = 8'h00;
    mem[16'h1BD9] = 8'h08; // POP RAX
    mem[16'h1BDA] = 8'h00;
    mem[16'h1BDB] = 8'h81; // ADDN RSP 8
    mem[16'h1BDC] = 8'h06;
    mem[16'h1BDD] = 8'h08;
    mem[16'h1BDE] = 8'h00;
    mem[16'h1BDF] = 8'h00;
    mem[16'h1BE0] = 8'h00;
    mem[16'h1BE1] = 8'h80; // ADD RAX RDI
    mem[16'h1BE2] = 8'h00;
    mem[16'h1BE3] = 8'h01;
    mem[16'h1BE4] = 8'h85; // SUBN RSP 8
    mem[16'h1BE5] = 8'h06;
    mem[16'h1BE6] = 8'h08;
    mem[16'h1BE7] = 8'h00;
    mem[16'h1BE8] = 8'h00;
    mem[16'h1BE9] = 8'h00;
    mem[16'h1BEA] = 8'h04; // PUSH RAX
    mem[16'h1BEB] = 8'h00;
    mem[16'h1BEC] = 8'h08; // POP RDI
    mem[16'h1BED] = 8'h01;
    mem[16'h1BEE] = 8'h81; // ADDN RSP 8
    mem[16'h1BEF] = 8'h06;
    mem[16'h1BF0] = 8'h08;
    mem[16'h1BF1] = 8'h00;
    mem[16'h1BF2] = 8'h00;
    mem[16'h1BF3] = 8'h00;
    mem[16'h1BF4] = 8'h08; // POP RAX
    mem[16'h1BF5] = 8'h00;
    mem[16'h1BF6] = 8'h81; // ADDN RSP 8
    mem[16'h1BF7] = 8'h06;
    mem[16'h1BF8] = 8'h08;
    mem[16'h1BF9] = 8'h00;
    mem[16'h1BFA] = 8'h00;
    mem[16'h1BFB] = 8'h00;
    mem[16'h1BFC] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h1BFD] = 8'h00;
    mem[16'h1BFE] = 8'h01;
    mem[16'h1BFF] = 8'h85; // SUBN RSP 8
    mem[16'h1C00] = 8'h06;
    mem[16'h1C01] = 8'h08;
    mem[16'h1C02] = 8'h00;
    mem[16'h1C03] = 8'h00;
    mem[16'h1C04] = 8'h00;
    mem[16'h1C05] = 8'h04; // PUSH RDI
    mem[16'h1C06] = 8'h01;
    mem[16'h1C07] = 8'h81; // ADDN RSP 8
    mem[16'h1C08] = 8'h06;
    mem[16'h1C09] = 8'h08;
    mem[16'h1C0A] = 8'h00;
    mem[16'h1C0B] = 8'h00;
    mem[16'h1C0C] = 8'h00;
    mem[16'h1C0D] = 8'h22; // JMP .Lbegin15
    mem[16'h1C0E] = 8'hA1;
    mem[16'h1C0F] = 8'h17;
    mem[16'h1C10] = 8'h00;
    mem[16'h1C11] = 8'h00;
    mem[16'h1C12] = 8'h00;
    mem[16'h1C13] = 8'h00;
    mem[16'h1C14] = 8'h00;
    mem[16'h1C15] = 8'h00;
                          // .Lend15:
    mem[16'h1C16] = 8'h40; // MOV RAX RBP
    mem[16'h1C17] = 8'h00;
    mem[16'h1C18] = 8'h05;
    mem[16'h1C19] = 8'h85; // SUBN RAX 4
    mem[16'h1C1A] = 8'h00;
    mem[16'h1C1B] = 8'h04;
    mem[16'h1C1C] = 8'h00;
    mem[16'h1C1D] = 8'h00;
    mem[16'h1C1E] = 8'h00;
    mem[16'h1C1F] = 8'h85; // SUBN RSP 8
    mem[16'h1C20] = 8'h06;
    mem[16'h1C21] = 8'h08;
    mem[16'h1C22] = 8'h00;
    mem[16'h1C23] = 8'h00;
    mem[16'h1C24] = 8'h00;
    mem[16'h1C25] = 8'h04; // PUSH RAX
    mem[16'h1C26] = 8'h00;
    mem[16'h1C27] = 8'h40; // MOV RAX RBP
    mem[16'h1C28] = 8'h00;
    mem[16'h1C29] = 8'h05;
    mem[16'h1C2A] = 8'h85; // SUBN RAX 4
    mem[16'h1C2B] = 8'h00;
    mem[16'h1C2C] = 8'h04;
    mem[16'h1C2D] = 8'h00;
    mem[16'h1C2E] = 8'h00;
    mem[16'h1C2F] = 8'h00;
    mem[16'h1C30] = 8'h85; // SUBN RSP 8
    mem[16'h1C31] = 8'h06;
    mem[16'h1C32] = 8'h08;
    mem[16'h1C33] = 8'h00;
    mem[16'h1C34] = 8'h00;
    mem[16'h1C35] = 8'h00;
    mem[16'h1C36] = 8'h04; // PUSH RAX
    mem[16'h1C37] = 8'h00;
    mem[16'h1C38] = 8'h08; // POP RAX
    mem[16'h1C39] = 8'h00;
    mem[16'h1C3A] = 8'h81; // ADDN RSP 8
    mem[16'h1C3B] = 8'h06;
    mem[16'h1C3C] = 8'h08;
    mem[16'h1C3D] = 8'h00;
    mem[16'h1C3E] = 8'h00;
    mem[16'h1C3F] = 8'h00;
    mem[16'h1C40] = 8'h48; // MOVRA4 RAX RAX
    mem[16'h1C41] = 8'h00;
    mem[16'h1C42] = 8'h00;
    mem[16'h1C43] = 8'h85; // SUBN RSP 8
    mem[16'h1C44] = 8'h06;
    mem[16'h1C45] = 8'h08;
    mem[16'h1C46] = 8'h00;
    mem[16'h1C47] = 8'h00;
    mem[16'h1C48] = 8'h00;
    mem[16'h1C49] = 8'h04; // PUSH RAX
    mem[16'h1C4A] = 8'h00;
    mem[16'h1C4B] = 8'h85; // SUBN RSP 8
    mem[16'h1C4C] = 8'h06;
    mem[16'h1C4D] = 8'h08;
    mem[16'h1C4E] = 8'h00;
    mem[16'h1C4F] = 8'h00;
    mem[16'h1C50] = 8'h00;
    mem[16'h1C51] = 8'h05; // PUSHN 1
    mem[16'h1C52] = 8'h00;
    mem[16'h1C53] = 8'h01;
    mem[16'h1C54] = 8'h00;
    mem[16'h1C55] = 8'h00;
    mem[16'h1C56] = 8'h00;
    mem[16'h1C57] = 8'h08; // POP RDI
    mem[16'h1C58] = 8'h01;
    mem[16'h1C59] = 8'h81; // ADDN RSP 8
    mem[16'h1C5A] = 8'h06;
    mem[16'h1C5B] = 8'h08;
    mem[16'h1C5C] = 8'h00;
    mem[16'h1C5D] = 8'h00;
    mem[16'h1C5E] = 8'h00;
    mem[16'h1C5F] = 8'h08; // POP RAX
    mem[16'h1C60] = 8'h00;
    mem[16'h1C61] = 8'h81; // ADDN RSP 8
    mem[16'h1C62] = 8'h06;
    mem[16'h1C63] = 8'h08;
    mem[16'h1C64] = 8'h00;
    mem[16'h1C65] = 8'h00;
    mem[16'h1C66] = 8'h00;
    mem[16'h1C67] = 8'h80; // ADD RAX RDI
    mem[16'h1C68] = 8'h00;
    mem[16'h1C69] = 8'h01;
    mem[16'h1C6A] = 8'h85; // SUBN RSP 8
    mem[16'h1C6B] = 8'h06;
    mem[16'h1C6C] = 8'h08;
    mem[16'h1C6D] = 8'h00;
    mem[16'h1C6E] = 8'h00;
    mem[16'h1C6F] = 8'h00;
    mem[16'h1C70] = 8'h04; // PUSH RAX
    mem[16'h1C71] = 8'h00;
    mem[16'h1C72] = 8'h08; // POP RDI
    mem[16'h1C73] = 8'h01;
    mem[16'h1C74] = 8'h81; // ADDN RSP 8
    mem[16'h1C75] = 8'h06;
    mem[16'h1C76] = 8'h08;
    mem[16'h1C77] = 8'h00;
    mem[16'h1C78] = 8'h00;
    mem[16'h1C79] = 8'h00;
    mem[16'h1C7A] = 8'h08; // POP RAX
    mem[16'h1C7B] = 8'h00;
    mem[16'h1C7C] = 8'h81; // ADDN RSP 8
    mem[16'h1C7D] = 8'h06;
    mem[16'h1C7E] = 8'h08;
    mem[16'h1C7F] = 8'h00;
    mem[16'h1C80] = 8'h00;
    mem[16'h1C81] = 8'h00;
    mem[16'h1C82] = 8'h58; // MOVAR4 RAX RDI
    mem[16'h1C83] = 8'h00;
    mem[16'h1C84] = 8'h01;
    mem[16'h1C85] = 8'h85; // SUBN RSP 8
    mem[16'h1C86] = 8'h06;
    mem[16'h1C87] = 8'h08;
    mem[16'h1C88] = 8'h00;
    mem[16'h1C89] = 8'h00;
    mem[16'h1C8A] = 8'h00;
    mem[16'h1C8B] = 8'h04; // PUSH RDI
    mem[16'h1C8C] = 8'h01;
    mem[16'h1C8D] = 8'h81; // ADDN RSP 8
    mem[16'h1C8E] = 8'h06;
    mem[16'h1C8F] = 8'h08;
    mem[16'h1C90] = 8'h00;
    mem[16'h1C91] = 8'h00;
    mem[16'h1C92] = 8'h00;
    mem[16'h1C93] = 8'h22; // JMP .Lbegin14
    mem[16'h1C94] = 8'hFC;
    mem[16'h1C95] = 8'h16;
    mem[16'h1C96] = 8'h00;
    mem[16'h1C97] = 8'h00;
    mem[16'h1C98] = 8'h00;
    mem[16'h1C99] = 8'h00;
    mem[16'h1C9A] = 8'h00;
    mem[16'h1C9B] = 8'h00;
                          // .Lend14:
    mem[16'h1C9C] = 8'h85; // SUBN RSP 8
    mem[16'h1C9D] = 8'h06;
    mem[16'h1C9E] = 8'h08;
    mem[16'h1C9F] = 8'h00;
    mem[16'h1CA0] = 8'h00;
    mem[16'h1CA1] = 8'h00;
    mem[16'h1CA2] = 8'h05; // PUSHN 0
    mem[16'h1CA3] = 8'h00;
    mem[16'h1CA4] = 8'h00;
    mem[16'h1CA5] = 8'h00;
    mem[16'h1CA6] = 8'h00;
    mem[16'h1CA7] = 8'h00;
    mem[16'h1CA8] = 8'h08; // POP RAX
    mem[16'h1CA9] = 8'h00;
    mem[16'h1CAA] = 8'h81; // ADDN RSP 8
    mem[16'h1CAB] = 8'h06;
    mem[16'h1CAC] = 8'h08;
    mem[16'h1CAD] = 8'h00;
    mem[16'h1CAE] = 8'h00;
    mem[16'h1CAF] = 8'h00;
    mem[16'h1CB0] = 8'h22; // JMP .Lreturn.eightqueen
    mem[16'h1CB1] = 8'hB9;
    mem[16'h1CB2] = 8'h1C;
    mem[16'h1CB3] = 8'h00;
    mem[16'h1CB4] = 8'h00;
    mem[16'h1CB5] = 8'h00;
    mem[16'h1CB6] = 8'h00;
    mem[16'h1CB7] = 8'h00;
    mem[16'h1CB8] = 8'h00;
                          // .Lreturn.eightqueen:
    mem[16'h1CB9] = 8'h40; // MOV RSP RBP
    mem[16'h1CBA] = 8'h06;
    mem[16'h1CBB] = 8'h05;
    mem[16'h1CBC] = 8'h08; // POP RBP
    mem[16'h1CBD] = 8'h05;
    mem[16'h1CBE] = 8'h81; // ADDN RSP 8
    mem[16'h1CBF] = 8'h06;
    mem[16'h1CC0] = 8'h08;
    mem[16'h1CC1] = 8'h00;
    mem[16'h1CC2] = 8'h00;
    mem[16'h1CC3] = 8'h00;
    mem[16'h1CC4] = 8'h08; // POP RBX
    mem[16'h1CC5] = 8'h07;
    mem[16'h1CC6] = 8'h81; // ADDN RSP 8
    mem[16'h1CC7] = 8'h06;
    mem[16'h1CC8] = 8'h08;
    mem[16'h1CC9] = 8'h00;
    mem[16'h1CCA] = 8'h00;
    mem[16'h1CCB] = 8'h00;
    mem[16'h1CCC] = 8'h20; // JMPR RBX
    mem[16'h1CCD] = 8'h07;
                          // main:
    mem[16'h1CCE] = 8'h85; // SUBN RSP 8
    mem[16'h1CCF] = 8'h06;
    mem[16'h1CD0] = 8'h08;
    mem[16'h1CD1] = 8'h00;
    mem[16'h1CD2] = 8'h00;
    mem[16'h1CD3] = 8'h00;
    mem[16'h1CD4] = 8'h04; // PUSH RBP
    mem[16'h1CD5] = 8'h05;
    mem[16'h1CD6] = 8'h40; // MOV RBP RSP
    mem[16'h1CD7] = 8'h05;
    mem[16'h1CD8] = 8'h06;
    mem[16'h1CD9] = 8'h85; // SUBN RSP 0
    mem[16'h1CDA] = 8'h06;
    mem[16'h1CDB] = 8'h00;
    mem[16'h1CDC] = 8'h00;
    mem[16'h1CDD] = 8'h00;
    mem[16'h1CDE] = 8'h00;
    mem[16'h1CDF] = 8'h85; // SUBN RSP 8
    mem[16'h1CE0] = 8'h06;
    mem[16'h1CE1] = 8'h08;
    mem[16'h1CE2] = 8'h00;
    mem[16'h1CE3] = 8'h00;
    mem[16'h1CE4] = 8'h00;
    mem[16'h1CE5] = 8'h05; // PUSHN 0
    mem[16'h1CE6] = 8'h00;
    mem[16'h1CE7] = 8'h00;
    mem[16'h1CE8] = 8'h00;
    mem[16'h1CE9] = 8'h00;
    mem[16'h1CEA] = 8'h00;
    mem[16'h1CEB] = 8'h08; // POP RDI
    mem[16'h1CEC] = 8'h01;
    mem[16'h1CED] = 8'h81; // ADDN RSP 8
    mem[16'h1CEE] = 8'h06;
    mem[16'h1CEF] = 8'h08;
    mem[16'h1CF0] = 8'h00;
    mem[16'h1CF1] = 8'h00;
    mem[16'h1CF2] = 8'h00;
    mem[16'h1CF3] = 8'h40; // MOV RAX RSP
    mem[16'h1CF4] = 8'h00;
    mem[16'h1CF5] = 8'h06;
    mem[16'h1CF6] = 8'h8D; // ANDN RAX 15
    mem[16'h1CF7] = 8'h00;
    mem[16'h1CF8] = 8'h0F;
    mem[16'h1CF9] = 8'h00;
    mem[16'h1CFA] = 8'h00;
    mem[16'h1CFB] = 8'h00;
    mem[16'h1CFC] = 8'h2A; // JNZ .Lcall20
    mem[16'h1CFD] = 8'h2D;
    mem[16'h1CFE] = 8'h1D;
    mem[16'h1CFF] = 8'h00;
    mem[16'h1D00] = 8'h00;
    mem[16'h1D01] = 8'h00;
    mem[16'h1D02] = 8'h00;
    mem[16'h1D03] = 8'h00;
    mem[16'h1D04] = 8'h00;
    mem[16'h1D05] = 8'h41; // MOVRN RAX 0
    mem[16'h1D06] = 8'h00;
    mem[16'h1D07] = 8'h00;
    mem[16'h1D08] = 8'h00;
    mem[16'h1D09] = 8'h00;
    mem[16'h1D0A] = 8'h00;
    mem[16'h1D0B] = 8'h0C; // MOVPC RBX
    mem[16'h1D0C] = 8'h07;
    mem[16'h1D0D] = 8'h81; // ADDN RBX 23
    mem[16'h1D0E] = 8'h07;
    mem[16'h1D0F] = 8'h17;
    mem[16'h1D10] = 8'h00;
    mem[16'h1D11] = 8'h00;
    mem[16'h1D12] = 8'h00;
    mem[16'h1D13] = 8'h85; // SUBN RSP 8
    mem[16'h1D14] = 8'h06;
    mem[16'h1D15] = 8'h08;
    mem[16'h1D16] = 8'h00;
    mem[16'h1D17] = 8'h00;
    mem[16'h1D18] = 8'h00;
    mem[16'h1D19] = 8'h04; // PUSH RBX
    mem[16'h1D1A] = 8'h07;
    mem[16'h1D1B] = 8'h22; // JMP eightqueen
    mem[16'h1D1C] = 8'h1D;
    mem[16'h1D1D] = 8'h16;
    mem[16'h1D1E] = 8'h00;
    mem[16'h1D1F] = 8'h00;
    mem[16'h1D20] = 8'h00;
    mem[16'h1D21] = 8'h00;
    mem[16'h1D22] = 8'h00;
    mem[16'h1D23] = 8'h00;
    mem[16'h1D24] = 8'h22; // JMP .Lend20
    mem[16'h1D25] = 8'h58;
    mem[16'h1D26] = 8'h1D;
    mem[16'h1D27] = 8'h00;
    mem[16'h1D28] = 8'h00;
    mem[16'h1D29] = 8'h00;
    mem[16'h1D2A] = 8'h00;
    mem[16'h1D2B] = 8'h00;
    mem[16'h1D2C] = 8'h00;
                          // .Lcall20:
    mem[16'h1D2D] = 8'h85; // SUBN RSP 8
    mem[16'h1D2E] = 8'h06;
    mem[16'h1D2F] = 8'h08;
    mem[16'h1D30] = 8'h00;
    mem[16'h1D31] = 8'h00;
    mem[16'h1D32] = 8'h00;
    mem[16'h1D33] = 8'h41; // MOVRN RAX 0
    mem[16'h1D34] = 8'h00;
    mem[16'h1D35] = 8'h00;
    mem[16'h1D36] = 8'h00;
    mem[16'h1D37] = 8'h00;
    mem[16'h1D38] = 8'h00;
    mem[16'h1D39] = 8'h0C; // MOVPC RBX
    mem[16'h1D3A] = 8'h07;
    mem[16'h1D3B] = 8'h81; // ADDN RBX 23
    mem[16'h1D3C] = 8'h07;
    mem[16'h1D3D] = 8'h17;
    mem[16'h1D3E] = 8'h00;
    mem[16'h1D3F] = 8'h00;
    mem[16'h1D40] = 8'h00;
    mem[16'h1D41] = 8'h85; // SUBN RSP 8
    mem[16'h1D42] = 8'h06;
    mem[16'h1D43] = 8'h08;
    mem[16'h1D44] = 8'h00;
    mem[16'h1D45] = 8'h00;
    mem[16'h1D46] = 8'h00;
    mem[16'h1D47] = 8'h04; // PUSH RBX
    mem[16'h1D48] = 8'h07;
    mem[16'h1D49] = 8'h22; // JMP eightqueen
    mem[16'h1D4A] = 8'h1D;
    mem[16'h1D4B] = 8'h16;
    mem[16'h1D4C] = 8'h00;
    mem[16'h1D4D] = 8'h00;
    mem[16'h1D4E] = 8'h00;
    mem[16'h1D4F] = 8'h00;
    mem[16'h1D50] = 8'h00;
    mem[16'h1D51] = 8'h00;
    mem[16'h1D52] = 8'h81; // ADDN RSP 8
    mem[16'h1D53] = 8'h06;
    mem[16'h1D54] = 8'h08;
    mem[16'h1D55] = 8'h00;
    mem[16'h1D56] = 8'h00;
    mem[16'h1D57] = 8'h00;
                          // .Lend20:
    mem[16'h1D58] = 8'h85; // SUBN RSP 8
    mem[16'h1D59] = 8'h06;
    mem[16'h1D5A] = 8'h08;
    mem[16'h1D5B] = 8'h00;
    mem[16'h1D5C] = 8'h00;
    mem[16'h1D5D] = 8'h00;
    mem[16'h1D5E] = 8'h04; // PUSH RAX
    mem[16'h1D5F] = 8'h00;
    mem[16'h1D60] = 8'h81; // ADDN RSP 8
    mem[16'h1D61] = 8'h06;
    mem[16'h1D62] = 8'h08;
    mem[16'h1D63] = 8'h00;
    mem[16'h1D64] = 8'h00;
    mem[16'h1D65] = 8'h00;
    mem[16'h1D66] = 8'h85; // SUBN RSP 8
    mem[16'h1D67] = 8'h06;
    mem[16'h1D68] = 8'h08;
    mem[16'h1D69] = 8'h00;
    mem[16'h1D6A] = 8'h00;
    mem[16'h1D6B] = 8'h00;
    mem[16'h1D6C] = 8'h05; // PUSHN 0
    mem[16'h1D6D] = 8'h00;
    mem[16'h1D6E] = 8'h00;
    mem[16'h1D6F] = 8'h00;
    mem[16'h1D70] = 8'h00;
    mem[16'h1D71] = 8'h00;
    mem[16'h1D72] = 8'h08; // POP RAX
    mem[16'h1D73] = 8'h00;
    mem[16'h1D74] = 8'h81; // ADDN RSP 8
    mem[16'h1D75] = 8'h06;
    mem[16'h1D76] = 8'h08;
    mem[16'h1D77] = 8'h00;
    mem[16'h1D78] = 8'h00;
    mem[16'h1D79] = 8'h00;
    mem[16'h1D7A] = 8'h22; // JMP .Lreturn.main
    mem[16'h1D7B] = 8'h83;
    mem[16'h1D7C] = 8'h1D;
    mem[16'h1D7D] = 8'h00;
    mem[16'h1D7E] = 8'h00;
    mem[16'h1D7F] = 8'h00;
    mem[16'h1D80] = 8'h00;
    mem[16'h1D81] = 8'h00;
    mem[16'h1D82] = 8'h00;
                          // .Lreturn.main:
    mem[16'h1D83] = 8'h00; // HLT
    mem[16'h1D84] = 8'h00;
    mem[16'h1D85] = 8'h40; // MOV RSP RBP
    mem[16'h1D86] = 8'h06;
    mem[16'h1D87] = 8'h05;
    mem[16'h1D88] = 8'h08; // POP RBP
    mem[16'h1D89] = 8'h05;
    mem[16'h1D8A] = 8'h81; // ADDN RSP 8
    mem[16'h1D8B] = 8'h06;
    mem[16'h1D8C] = 8'h08;
    mem[16'h1D8D] = 8'h00;
    mem[16'h1D8E] = 8'h00;
    mem[16'h1D8F] = 8'h00;
    mem[16'h1D90] = 8'h08; // POP RBX
    mem[16'h1D91] = 8'h07;
    mem[16'h1D92] = 8'h81; // ADDN RSP 8
    mem[16'h1D93] = 8'h06;
    mem[16'h1D94] = 8'h08;
    mem[16'h1D95] = 8'h00;
    mem[16'h1D96] = 8'h00;
    mem[16'h1D97] = 8'h00;
    mem[16'h1D98] = 8'h20; // JMPR RBX
    mem[16'h1D99] = 8'h07;
  end  
  
endmodule